magic
tech sky130A
timestamp 1650474576
<< nwell >>
rect -1600 0 -300 800
<< nmos >>
rect -1500 -600 -1400 -500
rect -700 -600 -600 -500
<< pmos >>
rect -1501 400 -1300 500
rect -800 200 -600 300
<< ndiff >>
rect -1500 -322 -1400 -300
rect -1500 -368 -1475 -322
rect -1417 -368 -1400 -322
rect -1500 -500 -1400 -368
rect -1000 -531 -700 -500
rect -1000 -571 -972 -531
rect -919 -571 -700 -531
rect -1000 -600 -700 -571
rect -600 -529 -400 -500
rect -600 -578 -474 -529
rect -417 -578 -400 -529
rect -600 -600 -400 -578
rect -1500 -927 -1400 -600
rect -1500 -981 -1474 -927
rect -1418 -981 -1400 -927
rect -1500 -1000 -1400 -981
<< pdiff >>
rect -1500 664 -1300 700
rect -1500 634 -1464 664
rect -1420 634 -1300 664
rect -1500 577 -1300 634
rect -1501 500 -1300 577
rect -1501 306 -1300 400
rect -1500 267 -1300 306
rect -1500 230 -1470 267
rect -1414 230 -1300 267
rect -1500 100 -1300 230
rect -1000 269 -800 300
rect -1000 235 -975 269
rect -932 235 -800 269
rect -1000 200 -800 235
rect -600 265 -400 300
rect -600 237 -467 265
rect -426 237 -400 265
rect -600 200 -400 237
<< ndiffc >>
rect -1475 -368 -1417 -322
rect -972 -571 -919 -531
rect -474 -578 -417 -529
rect -1474 -981 -1418 -927
<< pdiffc >>
rect -1464 634 -1420 664
rect -1470 230 -1414 267
rect -975 235 -932 269
rect -467 237 -426 265
<< poly >>
rect -1900 400 -1501 500
rect -1300 400 -1200 500
rect -1900 298 -1800 400
rect -1905 200 -1800 298
rect -1900 -238 -1800 200
rect -800 300 -600 400
rect -800 100 -600 200
rect -700 -124 -600 100
rect -700 -177 -675 -124
rect -616 -177 -600 -124
rect -700 -200 -600 -177
rect -1900 -263 -1874 -238
rect -1814 -263 -1800 -238
rect -1900 -500 -1800 -263
rect -700 -500 -600 -400
rect -1900 -600 -1500 -500
rect -1400 -600 -1300 -500
rect -700 -725 -600 -600
rect -700 -758 -676 -725
rect -614 -758 -600 -725
rect -700 -800 -600 -758
<< polycont >>
rect -675 -177 -616 -124
rect -1874 -263 -1814 -238
rect -676 -758 -614 -725
<< locali >>
rect -1481 664 -1412 679
rect -1481 634 -1464 664
rect -1420 634 -1412 664
rect -1481 623 -1412 634
rect -1486 267 -1407 276
rect -1486 230 -1470 267
rect -1414 230 -1407 267
rect -1486 222 -1407 230
rect -984 269 -917 274
rect -984 235 -975 269
rect -932 235 -917 269
rect -984 219 -917 235
rect -485 265 -413 278
rect -485 237 -467 265
rect -426 237 -413 265
rect -485 219 -413 237
rect -1388 -183 -1309 -113
rect -890 -190 -807 -110
rect -688 -124 -610 -112
rect -688 -177 -675 -124
rect -616 -177 -610 -124
rect -688 -187 -610 -177
rect -1890 -238 -1806 -227
rect -1890 -263 -1874 -238
rect -1814 -263 -1806 -238
rect -1890 -277 -1806 -263
rect -1492 -322 -1413 -307
rect -1492 -368 -1475 -322
rect -1417 -368 -1413 -322
rect -1492 -380 -1413 -368
rect -992 -531 -907 -516
rect -992 -571 -972 -531
rect -919 -571 -907 -531
rect -992 -584 -907 -571
rect -486 -529 -411 -515
rect -486 -578 -474 -529
rect -417 -578 -411 -529
rect -486 -586 -411 -578
rect -691 -725 -608 -711
rect -691 -758 -676 -725
rect -614 -758 -608 -725
rect -691 -776 -608 -758
rect -1494 -927 -1401 -913
rect -1494 -981 -1474 -927
rect -1418 -981 -1401 -927
rect -1494 -993 -1401 -981
<< metal1 >>
rect -1602 598 -209 781
rect -2600 200 -900 300
rect -500 200 -200 300
rect -1500 -100 -1400 200
rect -1500 -129 -1300 -100
rect -1500 -168 -1372 -129
rect -1317 -168 -1300 -129
rect -1500 -200 -1300 -168
rect -2600 -300 -1800 -200
rect -2400 -700 -2300 -300
rect -1500 -400 -1400 -200
rect -1200 -500 -1100 200
rect -300 -100 -200 200
rect -900 -127 -600 -100
rect -900 -179 -874 -127
rect -810 -179 -600 -127
rect -900 -200 -600 -179
rect -300 -200 100 -100
rect -300 -500 -200 -200
rect -1200 -600 -900 -500
rect -500 -600 -200 -500
rect -2400 -800 -600 -700
rect -1700 -922 -200 -900
rect -1704 -1110 -183 -922
<< via1 >>
rect -1372 -168 -1317 -129
rect -874 -179 -810 -127
<< metal2 >>
rect -1400 -127 -800 -100
rect -1400 -129 -874 -127
rect -1400 -168 -1372 -129
rect -1317 -168 -874 -129
rect -1400 -179 -874 -168
rect -810 -179 -800 -127
rect -1400 -200 -800 -179
<< labels >>
rlabel metal1 -1536 654 -1536 654 1 VDD!
rlabel metal1 -1600 -1100 -1600 -1100 5 GND!
rlabel metal1 -1655 -1058 -1655 -1058 5 GND!
rlabel metal1 -2554 266 -2554 266 5 Vin
rlabel metal1 -2558 -268 -2558 -268 5 S
rlabel metal1 61 -151 61 -151 5 Vout
<< end >>

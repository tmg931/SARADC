magic
tech sky130A
magscale 1 2
timestamp 1649880961
<< viali >>
rect 1501 11849 1535 11883
rect 6561 11849 6595 11883
rect 9229 11849 9263 11883
rect 10425 11849 10459 11883
rect 1685 11713 1719 11747
rect 2697 11713 2731 11747
rect 6377 11713 6411 11747
rect 7941 11713 7975 11747
rect 9413 11713 9447 11747
rect 10241 11713 10275 11747
rect 3801 11645 3835 11679
rect 4077 11577 4111 11611
rect 2881 11509 2915 11543
rect 4261 11509 4295 11543
rect 7757 11509 7791 11543
rect 10425 11237 10459 11271
rect 6929 11169 6963 11203
rect 8401 11169 8435 11203
rect 1777 11101 1811 11135
rect 5917 11101 5951 11135
rect 6653 11101 6687 11135
rect 10241 11101 10275 11135
rect 5641 11033 5675 11067
rect 4169 10965 4203 10999
rect 3709 10761 3743 10795
rect 9045 10761 9079 10795
rect 10149 10761 10183 10795
rect 7573 10693 7607 10727
rect 1777 10625 1811 10659
rect 6561 10625 6595 10659
rect 1409 10557 1443 10591
rect 5181 10557 5215 10591
rect 5457 10557 5491 10591
rect 7297 10557 7331 10591
rect 9873 10557 9907 10591
rect 10057 10557 10091 10591
rect 3203 10421 3237 10455
rect 6377 10421 6411 10455
rect 10517 10421 10551 10455
rect 1501 10217 1535 10251
rect 2697 10217 2731 10251
rect 4813 10217 4847 10251
rect 8953 10217 8987 10251
rect 10149 10217 10183 10251
rect 5549 10081 5583 10115
rect 9597 10081 9631 10115
rect 1685 10013 1719 10047
rect 2881 10013 2915 10047
rect 2973 10013 3007 10047
rect 3157 10013 3191 10047
rect 3249 10013 3283 10047
rect 4169 10013 4203 10047
rect 4353 10013 4387 10047
rect 4629 10013 4663 10047
rect 5273 10013 5307 10047
rect 7481 10013 7515 10047
rect 9321 10013 9355 10047
rect 10333 10013 10367 10047
rect 7665 9945 7699 9979
rect 7021 9877 7055 9911
rect 9413 9877 9447 9911
rect 3893 9673 3927 9707
rect 2145 9537 2179 9571
rect 4537 9537 4571 9571
rect 4813 9537 4847 9571
rect 4997 9537 5031 9571
rect 2421 9469 2455 9503
rect 8493 9469 8527 9503
rect 8769 9469 8803 9503
rect 10517 9469 10551 9503
rect 4353 9333 4387 9367
rect 4537 9129 4571 9163
rect 6929 8993 6963 9027
rect 2053 8925 2087 8959
rect 4721 8925 4755 8959
rect 4997 8925 5031 8959
rect 5181 8925 5215 8959
rect 6653 8925 6687 8959
rect 1869 8789 1903 8823
rect 8401 8789 8435 8823
rect 7021 8585 7055 8619
rect 9229 8585 9263 8619
rect 1685 8517 1719 8551
rect 4353 8517 4387 8551
rect 7757 8517 7791 8551
rect 1409 8449 1443 8483
rect 4077 8449 4111 8483
rect 6377 8449 6411 8483
rect 6561 8449 6595 8483
rect 6837 8449 6871 8483
rect 3157 8381 3191 8415
rect 7481 8381 7515 8415
rect 5825 8313 5859 8347
rect 2237 8041 2271 8075
rect 3801 8041 3835 8075
rect 8033 8041 8067 8075
rect 8953 8041 8987 8075
rect 2789 7905 2823 7939
rect 2605 7837 2639 7871
rect 5549 7837 5583 7871
rect 6285 7837 6319 7871
rect 9137 7837 9171 7871
rect 9413 7837 9447 7871
rect 9597 7837 9631 7871
rect 10241 7837 10275 7871
rect 5273 7769 5307 7803
rect 6561 7769 6595 7803
rect 2697 7701 2731 7735
rect 10425 7701 10459 7735
rect 4905 7497 4939 7531
rect 7941 7497 7975 7531
rect 2881 7429 2915 7463
rect 4445 7429 4479 7463
rect 3157 7361 3191 7395
rect 4537 7361 4571 7395
rect 7573 7361 7607 7395
rect 4261 7293 4295 7327
rect 7389 7293 7423 7327
rect 7481 7293 7515 7327
rect 10241 7293 10275 7327
rect 10517 7293 10551 7327
rect 8769 7225 8803 7259
rect 1409 7157 1443 7191
rect 1501 6885 1535 6919
rect 7297 6817 7331 6851
rect 1685 6749 1719 6783
rect 5549 6749 5583 6783
rect 9137 6749 9171 6783
rect 9321 6749 9355 6783
rect 9597 6749 9631 6783
rect 5825 6681 5859 6715
rect 9781 6613 9815 6647
rect 5825 6409 5859 6443
rect 6837 6409 6871 6443
rect 10149 6409 10183 6443
rect 2053 6341 2087 6375
rect 6929 6273 6963 6307
rect 1777 6205 1811 6239
rect 4077 6205 4111 6239
rect 4353 6205 4387 6239
rect 8401 6205 8435 6239
rect 8677 6205 8711 6239
rect 3525 6069 3559 6103
rect 3801 5729 3835 5763
rect 8125 5729 8159 5763
rect 9045 5729 9079 5763
rect 2513 5661 2547 5695
rect 2697 5661 2731 5695
rect 2973 5661 3007 5695
rect 3985 5661 4019 5695
rect 4261 5661 4295 5695
rect 4445 5661 4479 5695
rect 8401 5661 8435 5695
rect 9229 5661 9263 5695
rect 3157 5525 3191 5559
rect 6653 5525 6687 5559
rect 9321 5525 9355 5559
rect 9689 5525 9723 5559
rect 4629 5321 4663 5355
rect 8769 5321 8803 5355
rect 3157 5253 3191 5287
rect 7849 5253 7883 5287
rect 10241 5253 10275 5287
rect 2881 5185 2915 5219
rect 5365 5185 5399 5219
rect 5641 5185 5675 5219
rect 5825 5185 5859 5219
rect 10517 5185 10551 5219
rect 8125 5117 8159 5151
rect 5181 4981 5215 5015
rect 6377 4981 6411 5015
rect 1409 4777 1443 4811
rect 3801 4777 3835 4811
rect 6193 4777 6227 4811
rect 2881 4641 2915 4675
rect 4353 4641 4387 4675
rect 5549 4641 5583 4675
rect 9321 4641 9355 4675
rect 3157 4573 3191 4607
rect 5457 4573 5491 4607
rect 6377 4573 6411 4607
rect 6653 4573 6687 4607
rect 6837 4573 6871 4607
rect 7573 4573 7607 4607
rect 7849 4573 7883 4607
rect 8033 4573 8067 4607
rect 10517 4573 10551 4607
rect 4169 4505 4203 4539
rect 4261 4437 4295 4471
rect 4997 4437 5031 4471
rect 5365 4437 5399 4471
rect 7389 4437 7423 4471
rect 5089 4233 5123 4267
rect 5457 4233 5491 4267
rect 10517 4233 10551 4267
rect 1685 4097 1719 4131
rect 2145 4097 2179 4131
rect 4261 4097 4295 4131
rect 5549 4029 5583 4063
rect 5733 4029 5767 4063
rect 7849 4029 7883 4063
rect 8125 4029 8159 4063
rect 8769 4029 8803 4063
rect 9045 4029 9079 4063
rect 1501 3893 1535 3927
rect 2329 3893 2363 3927
rect 4077 3893 4111 3927
rect 6377 3893 6411 3927
rect 2605 3689 2639 3723
rect 5825 3689 5859 3723
rect 2053 3553 2087 3587
rect 2145 3553 2179 3587
rect 4077 3553 4111 3587
rect 4353 3553 4387 3587
rect 6929 3553 6963 3587
rect 9137 3553 9171 3587
rect 6653 3485 6687 3519
rect 9321 3485 9355 3519
rect 9597 3485 9631 3519
rect 9781 3485 9815 3519
rect 2237 3349 2271 3383
rect 8401 3349 8435 3383
rect 1409 3145 1443 3179
rect 5365 3145 5399 3179
rect 8953 3145 8987 3179
rect 2881 3077 2915 3111
rect 3893 3077 3927 3111
rect 7481 3077 7515 3111
rect 3157 3009 3191 3043
rect 3617 3009 3651 3043
rect 6469 3009 6503 3043
rect 7205 3009 7239 3043
rect 6653 2805 6687 2839
rect 8401 2601 8435 2635
rect 2053 2533 2087 2567
rect 4169 2465 4203 2499
rect 6653 2465 6687 2499
rect 6929 2465 6963 2499
rect 3801 2397 3835 2431
rect 9505 2397 9539 2431
rect 10241 2397 10275 2431
rect 1869 2329 1903 2363
rect 9689 2261 9723 2295
rect 10425 2261 10459 2295
<< metal1 >>
rect 1104 11994 11224 12016
rect 1104 11942 4323 11994
rect 4375 11942 4387 11994
rect 4439 11942 4451 11994
rect 4503 11942 4515 11994
rect 4567 11942 4579 11994
rect 4631 11942 7696 11994
rect 7748 11942 7760 11994
rect 7812 11942 7824 11994
rect 7876 11942 7888 11994
rect 7940 11942 7952 11994
rect 8004 11942 11224 11994
rect 1104 11920 11224 11942
rect 1486 11880 1492 11892
rect 1447 11852 1492 11880
rect 1486 11840 1492 11852
rect 1544 11840 1550 11892
rect 5810 11840 5816 11892
rect 5868 11880 5874 11892
rect 6549 11883 6607 11889
rect 6549 11880 6561 11883
rect 5868 11852 6561 11880
rect 5868 11840 5874 11852
rect 6549 11849 6561 11852
rect 6595 11849 6607 11883
rect 9214 11880 9220 11892
rect 9175 11852 9220 11880
rect 6549 11843 6607 11849
rect 9214 11840 9220 11852
rect 9272 11840 9278 11892
rect 10413 11883 10471 11889
rect 10413 11849 10425 11883
rect 10459 11880 10471 11883
rect 12250 11880 12256 11892
rect 10459 11852 12256 11880
rect 10459 11849 10471 11852
rect 10413 11843 10471 11849
rect 12250 11840 12256 11852
rect 12308 11840 12314 11892
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11744 1731 11747
rect 2498 11744 2504 11756
rect 1719 11716 2504 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 2498 11704 2504 11716
rect 2556 11704 2562 11756
rect 2682 11744 2688 11756
rect 2643 11716 2688 11744
rect 2682 11704 2688 11716
rect 2740 11704 2746 11756
rect 5718 11704 5724 11756
rect 5776 11744 5782 11756
rect 6365 11747 6423 11753
rect 6365 11744 6377 11747
rect 5776 11716 6377 11744
rect 5776 11704 5782 11716
rect 6365 11713 6377 11716
rect 6411 11713 6423 11747
rect 6365 11707 6423 11713
rect 7929 11747 7987 11753
rect 7929 11713 7941 11747
rect 7975 11744 7987 11747
rect 8938 11744 8944 11756
rect 7975 11716 8944 11744
rect 7975 11713 7987 11716
rect 7929 11707 7987 11713
rect 8938 11704 8944 11716
rect 8996 11704 9002 11756
rect 9030 11704 9036 11756
rect 9088 11744 9094 11756
rect 9401 11747 9459 11753
rect 9401 11744 9413 11747
rect 9088 11716 9413 11744
rect 9088 11704 9094 11716
rect 9401 11713 9413 11716
rect 9447 11713 9459 11747
rect 9401 11707 9459 11713
rect 10134 11704 10140 11756
rect 10192 11744 10198 11756
rect 10229 11747 10287 11753
rect 10229 11744 10241 11747
rect 10192 11716 10241 11744
rect 10192 11704 10198 11716
rect 10229 11713 10241 11716
rect 10275 11713 10287 11747
rect 10229 11707 10287 11713
rect 3789 11679 3847 11685
rect 3789 11676 3801 11679
rect 2976 11648 3801 11676
rect 2976 11552 3004 11648
rect 3789 11645 3801 11648
rect 3835 11645 3847 11679
rect 3789 11639 3847 11645
rect 3694 11568 3700 11620
rect 3752 11608 3758 11620
rect 4065 11611 4123 11617
rect 4065 11608 4077 11611
rect 3752 11580 4077 11608
rect 3752 11568 3758 11580
rect 4065 11577 4077 11580
rect 4111 11577 4123 11611
rect 4065 11571 4123 11577
rect 2869 11543 2927 11549
rect 2869 11509 2881 11543
rect 2915 11540 2927 11543
rect 2958 11540 2964 11552
rect 2915 11512 2964 11540
rect 2915 11509 2927 11512
rect 2869 11503 2927 11509
rect 2958 11500 2964 11512
rect 3016 11500 3022 11552
rect 4249 11543 4307 11549
rect 4249 11509 4261 11543
rect 4295 11540 4307 11543
rect 6546 11540 6552 11552
rect 4295 11512 6552 11540
rect 4295 11509 4307 11512
rect 4249 11503 4307 11509
rect 6546 11500 6552 11512
rect 6604 11500 6610 11552
rect 7558 11500 7564 11552
rect 7616 11540 7622 11552
rect 7745 11543 7803 11549
rect 7745 11540 7757 11543
rect 7616 11512 7757 11540
rect 7616 11500 7622 11512
rect 7745 11509 7757 11512
rect 7791 11509 7803 11543
rect 7745 11503 7803 11509
rect 1104 11450 11224 11472
rect 1104 11398 2636 11450
rect 2688 11398 2700 11450
rect 2752 11398 2764 11450
rect 2816 11398 2828 11450
rect 2880 11398 2892 11450
rect 2944 11398 6010 11450
rect 6062 11398 6074 11450
rect 6126 11398 6138 11450
rect 6190 11398 6202 11450
rect 6254 11398 6266 11450
rect 6318 11398 9383 11450
rect 9435 11398 9447 11450
rect 9499 11398 9511 11450
rect 9563 11398 9575 11450
rect 9627 11398 9639 11450
rect 9691 11398 11224 11450
rect 1104 11376 11224 11398
rect 10410 11268 10416 11280
rect 10371 11240 10416 11268
rect 10410 11228 10416 11240
rect 10468 11228 10474 11280
rect 6917 11203 6975 11209
rect 6917 11169 6929 11203
rect 6963 11200 6975 11203
rect 8389 11203 8447 11209
rect 6963 11172 8340 11200
rect 6963 11169 6975 11172
rect 6917 11163 6975 11169
rect 1762 11132 1768 11144
rect 1723 11104 1768 11132
rect 1762 11092 1768 11104
rect 1820 11092 1826 11144
rect 5902 11092 5908 11144
rect 5960 11132 5966 11144
rect 6641 11135 6699 11141
rect 6641 11132 6653 11135
rect 5960 11104 6653 11132
rect 5960 11092 5966 11104
rect 6641 11101 6653 11104
rect 6687 11101 6699 11135
rect 8312 11132 8340 11172
rect 8389 11169 8401 11203
rect 8435 11200 8447 11203
rect 10134 11200 10140 11212
rect 8435 11172 10140 11200
rect 8435 11169 8447 11172
rect 8389 11163 8447 11169
rect 10134 11160 10140 11172
rect 10192 11160 10198 11212
rect 10042 11132 10048 11144
rect 8312 11104 10048 11132
rect 6641 11095 6699 11101
rect 10042 11092 10048 11104
rect 10100 11092 10106 11144
rect 10226 11132 10232 11144
rect 10187 11104 10232 11132
rect 10226 11092 10232 11104
rect 10284 11092 10290 11144
rect 4062 11024 4068 11076
rect 4120 11064 4126 11076
rect 5626 11064 5632 11076
rect 4120 11036 4462 11064
rect 5587 11036 5632 11064
rect 4120 11024 4126 11036
rect 5626 11024 5632 11036
rect 5684 11024 5690 11076
rect 8662 11064 8668 11076
rect 8142 11036 8668 11064
rect 8662 11024 8668 11036
rect 8720 11024 8726 11076
rect 4154 10996 4160 11008
rect 4115 10968 4160 10996
rect 4154 10956 4160 10968
rect 4212 10956 4218 11008
rect 1104 10906 11224 10928
rect 1104 10854 4323 10906
rect 4375 10854 4387 10906
rect 4439 10854 4451 10906
rect 4503 10854 4515 10906
rect 4567 10854 4579 10906
rect 4631 10854 7696 10906
rect 7748 10854 7760 10906
rect 7812 10854 7824 10906
rect 7876 10854 7888 10906
rect 7940 10854 7952 10906
rect 8004 10854 11224 10906
rect 1104 10832 11224 10854
rect 3694 10792 3700 10804
rect 3655 10764 3700 10792
rect 3694 10752 3700 10764
rect 3752 10752 3758 10804
rect 9030 10792 9036 10804
rect 8991 10764 9036 10792
rect 9030 10752 9036 10764
rect 9088 10752 9094 10804
rect 10134 10792 10140 10804
rect 10095 10764 10140 10792
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 7558 10724 7564 10736
rect 1762 10656 1768 10668
rect 1723 10628 1768 10656
rect 1762 10616 1768 10628
rect 1820 10616 1826 10668
rect 2792 10656 2820 10710
rect 7519 10696 7564 10724
rect 7558 10684 7564 10696
rect 7616 10684 7622 10736
rect 3418 10656 3424 10668
rect 2792 10628 3424 10656
rect 3418 10616 3424 10628
rect 3476 10656 3482 10668
rect 4062 10656 4068 10668
rect 3476 10628 4068 10656
rect 3476 10616 3482 10628
rect 4062 10616 4068 10628
rect 4120 10616 4126 10668
rect 6546 10656 6552 10668
rect 6507 10628 6552 10656
rect 6546 10616 6552 10628
rect 6604 10616 6610 10668
rect 8662 10616 8668 10668
rect 8720 10616 8726 10668
rect 1394 10588 1400 10600
rect 1355 10560 1400 10588
rect 1394 10548 1400 10560
rect 1452 10548 1458 10600
rect 3050 10548 3056 10600
rect 3108 10588 3114 10600
rect 5169 10591 5227 10597
rect 5169 10588 5181 10591
rect 3108 10560 5181 10588
rect 3108 10548 3114 10560
rect 5169 10557 5181 10560
rect 5215 10557 5227 10591
rect 5169 10551 5227 10557
rect 5445 10591 5503 10597
rect 5445 10557 5457 10591
rect 5491 10588 5503 10591
rect 5810 10588 5816 10600
rect 5491 10560 5816 10588
rect 5491 10557 5503 10560
rect 5445 10551 5503 10557
rect 5810 10548 5816 10560
rect 5868 10588 5874 10600
rect 7285 10591 7343 10597
rect 7285 10588 7297 10591
rect 5868 10560 7297 10588
rect 5868 10548 5874 10560
rect 7285 10557 7297 10560
rect 7331 10557 7343 10591
rect 7285 10551 7343 10557
rect 9766 10548 9772 10600
rect 9824 10588 9830 10600
rect 9861 10591 9919 10597
rect 9861 10588 9873 10591
rect 9824 10560 9873 10588
rect 9824 10548 9830 10560
rect 9861 10557 9873 10560
rect 9907 10557 9919 10591
rect 9861 10551 9919 10557
rect 9950 10548 9956 10600
rect 10008 10588 10014 10600
rect 10045 10591 10103 10597
rect 10045 10588 10057 10591
rect 10008 10560 10057 10588
rect 10008 10548 10014 10560
rect 10045 10557 10057 10560
rect 10091 10557 10103 10591
rect 10045 10551 10103 10557
rect 3142 10412 3148 10464
rect 3200 10461 3206 10464
rect 3200 10455 3249 10461
rect 3200 10421 3203 10455
rect 3237 10421 3249 10455
rect 3200 10415 3249 10421
rect 3200 10412 3206 10415
rect 5534 10412 5540 10464
rect 5592 10452 5598 10464
rect 6365 10455 6423 10461
rect 6365 10452 6377 10455
rect 5592 10424 6377 10452
rect 5592 10412 5598 10424
rect 6365 10421 6377 10424
rect 6411 10421 6423 10455
rect 6365 10415 6423 10421
rect 10318 10412 10324 10464
rect 10376 10452 10382 10464
rect 10505 10455 10563 10461
rect 10505 10452 10517 10455
rect 10376 10424 10517 10452
rect 10376 10412 10382 10424
rect 10505 10421 10517 10424
rect 10551 10421 10563 10455
rect 10505 10415 10563 10421
rect 1104 10362 11224 10384
rect 1104 10310 2636 10362
rect 2688 10310 2700 10362
rect 2752 10310 2764 10362
rect 2816 10310 2828 10362
rect 2880 10310 2892 10362
rect 2944 10310 6010 10362
rect 6062 10310 6074 10362
rect 6126 10310 6138 10362
rect 6190 10310 6202 10362
rect 6254 10310 6266 10362
rect 6318 10310 9383 10362
rect 9435 10310 9447 10362
rect 9499 10310 9511 10362
rect 9563 10310 9575 10362
rect 9627 10310 9639 10362
rect 9691 10310 11224 10362
rect 1104 10288 11224 10310
rect 1486 10248 1492 10260
rect 1447 10220 1492 10248
rect 1486 10208 1492 10220
rect 1544 10208 1550 10260
rect 2685 10251 2743 10257
rect 2685 10217 2697 10251
rect 2731 10248 2743 10251
rect 3050 10248 3056 10260
rect 2731 10220 3056 10248
rect 2731 10217 2743 10220
rect 2685 10211 2743 10217
rect 3050 10208 3056 10220
rect 3108 10208 3114 10260
rect 4801 10251 4859 10257
rect 4801 10217 4813 10251
rect 4847 10248 4859 10251
rect 5626 10248 5632 10260
rect 4847 10220 5632 10248
rect 4847 10217 4859 10220
rect 4801 10211 4859 10217
rect 5626 10208 5632 10220
rect 5684 10208 5690 10260
rect 8938 10248 8944 10260
rect 8899 10220 8944 10248
rect 8938 10208 8944 10220
rect 8996 10208 9002 10260
rect 10042 10208 10048 10260
rect 10100 10248 10106 10260
rect 10137 10251 10195 10257
rect 10137 10248 10149 10251
rect 10100 10220 10149 10248
rect 10100 10208 10106 10220
rect 10137 10217 10149 10220
rect 10183 10217 10195 10251
rect 10137 10211 10195 10217
rect 4154 10180 4160 10192
rect 1688 10152 4160 10180
rect 1688 10053 1716 10152
rect 4154 10140 4160 10152
rect 4212 10180 4218 10192
rect 4212 10152 4384 10180
rect 4212 10140 4218 10152
rect 3694 10112 3700 10124
rect 2976 10084 3700 10112
rect 1673 10047 1731 10053
rect 1673 10013 1685 10047
rect 1719 10013 1731 10047
rect 2866 10044 2872 10056
rect 2827 10016 2872 10044
rect 1673 10007 1731 10013
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 2976 10053 3004 10084
rect 3694 10072 3700 10084
rect 3752 10072 3758 10124
rect 2961 10047 3019 10053
rect 2961 10013 2973 10047
rect 3007 10013 3019 10047
rect 3142 10044 3148 10056
rect 3103 10016 3148 10044
rect 2961 10007 3019 10013
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 3237 10047 3295 10053
rect 3237 10013 3249 10047
rect 3283 10044 3295 10047
rect 4154 10044 4160 10056
rect 3283 10016 3924 10044
rect 4115 10016 4160 10044
rect 3283 10013 3295 10016
rect 3237 10007 3295 10013
rect 3896 9988 3924 10016
rect 4154 10004 4160 10016
rect 4212 10004 4218 10056
rect 4356 10053 4384 10152
rect 5534 10112 5540 10124
rect 5495 10084 5540 10112
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 7006 10112 7012 10124
rect 6656 10084 7012 10112
rect 4341 10047 4399 10053
rect 4341 10013 4353 10047
rect 4387 10013 4399 10047
rect 4341 10007 4399 10013
rect 4617 10047 4675 10053
rect 4617 10013 4629 10047
rect 4663 10013 4675 10047
rect 4617 10007 4675 10013
rect 5261 10047 5319 10053
rect 5261 10013 5273 10047
rect 5307 10013 5319 10047
rect 6656 10030 6684 10084
rect 7006 10072 7012 10084
rect 7064 10072 7070 10124
rect 9585 10115 9643 10121
rect 9585 10081 9597 10115
rect 9631 10112 9643 10115
rect 9766 10112 9772 10124
rect 9631 10084 9772 10112
rect 9631 10081 9643 10084
rect 9585 10075 9643 10081
rect 9766 10072 9772 10084
rect 9824 10072 9830 10124
rect 5261 10007 5319 10013
rect 3878 9936 3884 9988
rect 3936 9976 3942 9988
rect 4632 9976 4660 10007
rect 3936 9948 4660 9976
rect 3936 9936 3942 9948
rect 5276 9908 5304 10007
rect 6822 10004 6828 10056
rect 6880 10044 6886 10056
rect 7469 10047 7527 10053
rect 7469 10044 7481 10047
rect 6880 10016 7481 10044
rect 6880 10004 6886 10016
rect 7469 10013 7481 10016
rect 7515 10013 7527 10047
rect 7469 10007 7527 10013
rect 9030 10004 9036 10056
rect 9088 10044 9094 10056
rect 9309 10047 9367 10053
rect 9309 10044 9321 10047
rect 9088 10016 9321 10044
rect 9088 10004 9094 10016
rect 9309 10013 9321 10016
rect 9355 10013 9367 10047
rect 10318 10044 10324 10056
rect 10279 10016 10324 10044
rect 9309 10007 9367 10013
rect 10318 10004 10324 10016
rect 10376 10004 10382 10056
rect 7653 9979 7711 9985
rect 7653 9976 7665 9979
rect 7024 9948 7665 9976
rect 5810 9908 5816 9920
rect 5276 9880 5816 9908
rect 5810 9868 5816 9880
rect 5868 9908 5874 9920
rect 6546 9908 6552 9920
rect 5868 9880 6552 9908
rect 5868 9868 5874 9880
rect 6546 9868 6552 9880
rect 6604 9868 6610 9920
rect 6914 9868 6920 9920
rect 6972 9908 6978 9920
rect 7024 9917 7052 9948
rect 7653 9945 7665 9948
rect 7699 9945 7711 9979
rect 7653 9939 7711 9945
rect 7009 9911 7067 9917
rect 7009 9908 7021 9911
rect 6972 9880 7021 9908
rect 6972 9868 6978 9880
rect 7009 9877 7021 9880
rect 7055 9877 7067 9911
rect 7009 9871 7067 9877
rect 8386 9868 8392 9920
rect 8444 9908 8450 9920
rect 9401 9911 9459 9917
rect 9401 9908 9413 9911
rect 8444 9880 9413 9908
rect 8444 9868 8450 9880
rect 9401 9877 9413 9880
rect 9447 9877 9459 9911
rect 9401 9871 9459 9877
rect 1104 9818 11224 9840
rect 1104 9766 4323 9818
rect 4375 9766 4387 9818
rect 4439 9766 4451 9818
rect 4503 9766 4515 9818
rect 4567 9766 4579 9818
rect 4631 9766 7696 9818
rect 7748 9766 7760 9818
rect 7812 9766 7824 9818
rect 7876 9766 7888 9818
rect 7940 9766 7952 9818
rect 8004 9766 11224 9818
rect 1104 9744 11224 9766
rect 3878 9704 3884 9716
rect 3839 9676 3884 9704
rect 3878 9664 3884 9676
rect 3936 9664 3942 9716
rect 4154 9664 4160 9716
rect 4212 9704 4218 9716
rect 6822 9704 6828 9716
rect 4212 9676 6828 9704
rect 4212 9664 4218 9676
rect 6822 9664 6828 9676
rect 6880 9664 6886 9716
rect 3418 9596 3424 9648
rect 3476 9596 3482 9648
rect 7006 9596 7012 9648
rect 7064 9636 7070 9648
rect 8202 9636 8208 9648
rect 7064 9608 8208 9636
rect 7064 9596 7070 9608
rect 8202 9596 8208 9608
rect 8260 9636 8266 9648
rect 8662 9636 8668 9648
rect 8260 9608 8668 9636
rect 8260 9596 8266 9608
rect 8662 9596 8668 9608
rect 8720 9636 8726 9648
rect 8720 9608 9246 9636
rect 8720 9596 8726 9608
rect 1394 9528 1400 9580
rect 1452 9568 1458 9580
rect 2133 9571 2191 9577
rect 2133 9568 2145 9571
rect 1452 9540 2145 9568
rect 1452 9528 1458 9540
rect 2133 9537 2145 9540
rect 2179 9537 2191 9571
rect 2133 9531 2191 9537
rect 4525 9571 4583 9577
rect 4525 9537 4537 9571
rect 4571 9537 4583 9571
rect 4798 9568 4804 9580
rect 4759 9540 4804 9568
rect 4525 9531 4583 9537
rect 2406 9500 2412 9512
rect 2319 9472 2412 9500
rect 2406 9460 2412 9472
rect 2464 9500 2470 9512
rect 4540 9500 4568 9531
rect 4798 9528 4804 9540
rect 4856 9528 4862 9580
rect 4985 9571 5043 9577
rect 4985 9537 4997 9571
rect 5031 9568 5043 9571
rect 5350 9568 5356 9580
rect 5031 9540 5356 9568
rect 5031 9537 5043 9540
rect 4985 9531 5043 9537
rect 5350 9528 5356 9540
rect 5408 9528 5414 9580
rect 4890 9500 4896 9512
rect 2464 9472 3556 9500
rect 4540 9472 4896 9500
rect 2464 9460 2470 9472
rect 3528 9432 3556 9472
rect 4890 9460 4896 9472
rect 4948 9460 4954 9512
rect 6638 9460 6644 9512
rect 6696 9500 6702 9512
rect 8481 9503 8539 9509
rect 8481 9500 8493 9503
rect 6696 9472 8493 9500
rect 6696 9460 6702 9472
rect 8481 9469 8493 9472
rect 8527 9469 8539 9503
rect 8481 9463 8539 9469
rect 8757 9503 8815 9509
rect 8757 9469 8769 9503
rect 8803 9500 8815 9503
rect 9214 9500 9220 9512
rect 8803 9472 9220 9500
rect 8803 9469 8815 9472
rect 8757 9463 8815 9469
rect 9214 9460 9220 9472
rect 9272 9460 9278 9512
rect 9766 9460 9772 9512
rect 9824 9500 9830 9512
rect 10505 9503 10563 9509
rect 10505 9500 10517 9503
rect 9824 9472 10517 9500
rect 9824 9460 9830 9472
rect 10505 9469 10517 9472
rect 10551 9469 10563 9503
rect 10505 9463 10563 9469
rect 3528 9404 6914 9432
rect 4246 9324 4252 9376
rect 4304 9364 4310 9376
rect 4341 9367 4399 9373
rect 4341 9364 4353 9367
rect 4304 9336 4353 9364
rect 4304 9324 4310 9336
rect 4341 9333 4353 9336
rect 4387 9333 4399 9367
rect 6886 9364 6914 9404
rect 9766 9364 9772 9376
rect 6886 9336 9772 9364
rect 4341 9327 4399 9333
rect 9766 9324 9772 9336
rect 9824 9324 9830 9376
rect 1104 9274 11224 9296
rect 1104 9222 2636 9274
rect 2688 9222 2700 9274
rect 2752 9222 2764 9274
rect 2816 9222 2828 9274
rect 2880 9222 2892 9274
rect 2944 9222 6010 9274
rect 6062 9222 6074 9274
rect 6126 9222 6138 9274
rect 6190 9222 6202 9274
rect 6254 9222 6266 9274
rect 6318 9222 9383 9274
rect 9435 9222 9447 9274
rect 9499 9222 9511 9274
rect 9563 9222 9575 9274
rect 9627 9222 9639 9274
rect 9691 9222 11224 9274
rect 1104 9200 11224 9222
rect 4525 9163 4583 9169
rect 4525 9129 4537 9163
rect 4571 9160 4583 9163
rect 4798 9160 4804 9172
rect 4571 9132 4804 9160
rect 4571 9129 4583 9132
rect 4525 9123 4583 9129
rect 4798 9120 4804 9132
rect 4856 9120 4862 9172
rect 4154 8984 4160 9036
rect 4212 9024 4218 9036
rect 6917 9027 6975 9033
rect 4212 8996 4844 9024
rect 4212 8984 4218 8996
rect 4816 8968 4844 8996
rect 6917 8993 6929 9027
rect 6963 9024 6975 9027
rect 8938 9024 8944 9036
rect 6963 8996 8944 9024
rect 6963 8993 6975 8996
rect 6917 8987 6975 8993
rect 8938 8984 8944 8996
rect 8996 8984 9002 9036
rect 2038 8956 2044 8968
rect 1999 8928 2044 8956
rect 2038 8916 2044 8928
rect 2096 8916 2102 8968
rect 4706 8956 4712 8968
rect 4667 8928 4712 8956
rect 4706 8916 4712 8928
rect 4764 8916 4770 8968
rect 4798 8916 4804 8968
rect 4856 8956 4862 8968
rect 4985 8959 5043 8965
rect 4985 8956 4997 8959
rect 4856 8928 4997 8956
rect 4856 8916 4862 8928
rect 4985 8925 4997 8928
rect 5031 8925 5043 8959
rect 4985 8919 5043 8925
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8956 5227 8959
rect 5258 8956 5264 8968
rect 5215 8928 5264 8956
rect 5215 8925 5227 8928
rect 5169 8919 5227 8925
rect 5258 8916 5264 8928
rect 5316 8916 5322 8968
rect 6638 8956 6644 8968
rect 6599 8928 6644 8956
rect 6638 8916 6644 8928
rect 6696 8916 6702 8968
rect 8202 8956 8208 8968
rect 8050 8928 8208 8956
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 10226 8888 10232 8900
rect 8220 8860 10232 8888
rect 1670 8780 1676 8832
rect 1728 8820 1734 8832
rect 1857 8823 1915 8829
rect 1857 8820 1869 8823
rect 1728 8792 1869 8820
rect 1728 8780 1734 8792
rect 1857 8789 1869 8792
rect 1903 8789 1915 8823
rect 1857 8783 1915 8789
rect 5350 8780 5356 8832
rect 5408 8820 5414 8832
rect 8220 8820 8248 8860
rect 10226 8848 10232 8860
rect 10284 8848 10290 8900
rect 8386 8820 8392 8832
rect 5408 8792 8248 8820
rect 8347 8792 8392 8820
rect 5408 8780 5414 8792
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 1104 8730 11224 8752
rect 1104 8678 4323 8730
rect 4375 8678 4387 8730
rect 4439 8678 4451 8730
rect 4503 8678 4515 8730
rect 4567 8678 4579 8730
rect 4631 8678 7696 8730
rect 7748 8678 7760 8730
rect 7812 8678 7824 8730
rect 7876 8678 7888 8730
rect 7940 8678 7952 8730
rect 8004 8678 11224 8730
rect 1104 8656 11224 8678
rect 1394 8576 1400 8628
rect 1452 8616 1458 8628
rect 3142 8616 3148 8628
rect 1452 8588 3148 8616
rect 1452 8576 1458 8588
rect 3142 8576 3148 8588
rect 3200 8616 3206 8628
rect 7009 8619 7067 8625
rect 3200 8588 4108 8616
rect 3200 8576 3206 8588
rect 1670 8548 1676 8560
rect 1631 8520 1676 8548
rect 1670 8508 1676 8520
rect 1728 8508 1734 8560
rect 3418 8548 3424 8560
rect 2898 8520 3424 8548
rect 3418 8508 3424 8520
rect 3476 8508 3482 8560
rect 1394 8480 1400 8492
rect 1355 8452 1400 8480
rect 1394 8440 1400 8452
rect 1452 8440 1458 8492
rect 2406 8372 2412 8424
rect 2464 8412 2470 8424
rect 3145 8415 3203 8421
rect 3145 8412 3157 8415
rect 2464 8384 3157 8412
rect 2464 8372 2470 8384
rect 3145 8381 3157 8384
rect 3191 8381 3203 8415
rect 3436 8412 3464 8508
rect 4080 8489 4108 8588
rect 7009 8585 7021 8619
rect 7055 8616 7067 8619
rect 8754 8616 8760 8628
rect 7055 8588 8760 8616
rect 7055 8585 7067 8588
rect 7009 8579 7067 8585
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 9214 8616 9220 8628
rect 9175 8588 9220 8616
rect 9214 8576 9220 8588
rect 9272 8576 9278 8628
rect 4246 8508 4252 8560
rect 4304 8548 4310 8560
rect 4341 8551 4399 8557
rect 4341 8548 4353 8551
rect 4304 8520 4353 8548
rect 4304 8508 4310 8520
rect 4341 8517 4353 8520
rect 4387 8517 4399 8551
rect 7374 8548 7380 8560
rect 4341 8511 4399 8517
rect 6840 8520 7380 8548
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8449 4123 8483
rect 6365 8483 6423 8489
rect 4065 8443 4123 8449
rect 3970 8412 3976 8424
rect 3436 8384 3976 8412
rect 3145 8375 3203 8381
rect 3970 8372 3976 8384
rect 4028 8412 4034 8424
rect 5460 8412 5488 8466
rect 6365 8449 6377 8483
rect 6411 8449 6423 8483
rect 6546 8480 6552 8492
rect 6507 8452 6552 8480
rect 6365 8443 6423 8449
rect 4028 8384 5488 8412
rect 6380 8412 6408 8443
rect 6546 8440 6552 8452
rect 6604 8440 6610 8492
rect 6840 8489 6868 8520
rect 7374 8508 7380 8520
rect 7432 8548 7438 8560
rect 7745 8551 7803 8557
rect 7745 8548 7757 8551
rect 7432 8520 7757 8548
rect 7432 8508 7438 8520
rect 7745 8517 7757 8520
rect 7791 8548 7803 8551
rect 8018 8548 8024 8560
rect 7791 8520 8024 8548
rect 7791 8517 7803 8520
rect 7745 8511 7803 8517
rect 8018 8508 8024 8520
rect 8076 8508 8082 8560
rect 8202 8508 8208 8560
rect 8260 8508 8266 8560
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8449 6883 8483
rect 6825 8443 6883 8449
rect 6914 8412 6920 8424
rect 6380 8384 6920 8412
rect 4028 8372 4034 8384
rect 6914 8372 6920 8384
rect 6972 8372 6978 8424
rect 7469 8415 7527 8421
rect 7469 8381 7481 8415
rect 7515 8381 7527 8415
rect 7469 8375 7527 8381
rect 5442 8304 5448 8356
rect 5500 8344 5506 8356
rect 5813 8347 5871 8353
rect 5813 8344 5825 8347
rect 5500 8316 5825 8344
rect 5500 8304 5506 8316
rect 5813 8313 5825 8316
rect 5859 8313 5871 8347
rect 5813 8307 5871 8313
rect 6638 8304 6644 8356
rect 6696 8344 6702 8356
rect 7484 8344 7512 8375
rect 6696 8316 7512 8344
rect 6696 8304 6702 8316
rect 1104 8186 11224 8208
rect 1104 8134 2636 8186
rect 2688 8134 2700 8186
rect 2752 8134 2764 8186
rect 2816 8134 2828 8186
rect 2880 8134 2892 8186
rect 2944 8134 6010 8186
rect 6062 8134 6074 8186
rect 6126 8134 6138 8186
rect 6190 8134 6202 8186
rect 6254 8134 6266 8186
rect 6318 8134 9383 8186
rect 9435 8134 9447 8186
rect 9499 8134 9511 8186
rect 9563 8134 9575 8186
rect 9627 8134 9639 8186
rect 9691 8134 11224 8186
rect 1104 8112 11224 8134
rect 2038 8032 2044 8084
rect 2096 8072 2102 8084
rect 2225 8075 2283 8081
rect 2225 8072 2237 8075
rect 2096 8044 2237 8072
rect 2096 8032 2102 8044
rect 2225 8041 2237 8044
rect 2271 8041 2283 8075
rect 2225 8035 2283 8041
rect 3789 8075 3847 8081
rect 3789 8041 3801 8075
rect 3835 8072 3847 8075
rect 4246 8072 4252 8084
rect 3835 8044 4252 8072
rect 3835 8041 3847 8044
rect 3789 8035 3847 8041
rect 4246 8032 4252 8044
rect 4304 8072 4310 8084
rect 4706 8072 4712 8084
rect 4304 8044 4712 8072
rect 4304 8032 4310 8044
rect 4706 8032 4712 8044
rect 4764 8032 4770 8084
rect 8018 8072 8024 8084
rect 7979 8044 8024 8072
rect 8018 8032 8024 8044
rect 8076 8032 8082 8084
rect 8938 8072 8944 8084
rect 8899 8044 8944 8072
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 8386 7964 8392 8016
rect 8444 8004 8450 8016
rect 8444 7976 9628 8004
rect 8444 7964 8450 7976
rect 2038 7896 2044 7948
rect 2096 7936 2102 7948
rect 2314 7936 2320 7948
rect 2096 7908 2320 7936
rect 2096 7896 2102 7908
rect 2314 7896 2320 7908
rect 2372 7936 2378 7948
rect 2777 7939 2835 7945
rect 2777 7936 2789 7939
rect 2372 7908 2789 7936
rect 2372 7896 2378 7908
rect 2777 7905 2789 7908
rect 2823 7905 2835 7939
rect 6638 7936 6644 7948
rect 2777 7899 2835 7905
rect 6288 7908 6644 7936
rect 2406 7828 2412 7880
rect 2464 7868 2470 7880
rect 2593 7871 2651 7877
rect 2593 7868 2605 7871
rect 2464 7840 2605 7868
rect 2464 7828 2470 7840
rect 2593 7837 2605 7840
rect 2639 7837 2651 7871
rect 2593 7831 2651 7837
rect 5534 7828 5540 7880
rect 5592 7868 5598 7880
rect 6288 7877 6316 7908
rect 6638 7896 6644 7908
rect 6696 7896 6702 7948
rect 8754 7896 8760 7948
rect 8812 7936 8818 7948
rect 8812 7908 9444 7936
rect 8812 7896 8818 7908
rect 6273 7871 6331 7877
rect 6273 7868 6285 7871
rect 5592 7840 6285 7868
rect 5592 7828 5598 7840
rect 6273 7837 6285 7840
rect 6319 7837 6331 7871
rect 6273 7831 6331 7837
rect 8018 7828 8024 7880
rect 8076 7868 8082 7880
rect 9416 7877 9444 7908
rect 9600 7877 9628 7976
rect 9125 7871 9183 7877
rect 9125 7868 9137 7871
rect 8076 7840 9137 7868
rect 8076 7828 8082 7840
rect 9125 7837 9137 7840
rect 9171 7837 9183 7871
rect 9125 7831 9183 7837
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 9585 7871 9643 7877
rect 9585 7837 9597 7871
rect 9631 7868 9643 7871
rect 10229 7871 10287 7877
rect 10229 7868 10241 7871
rect 9631 7840 10241 7868
rect 9631 7837 9643 7840
rect 9585 7831 9643 7837
rect 10229 7837 10241 7840
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 3970 7760 3976 7812
rect 4028 7800 4034 7812
rect 5258 7800 5264 7812
rect 4028 7772 4094 7800
rect 5219 7772 5264 7800
rect 4028 7760 4034 7772
rect 5258 7760 5264 7772
rect 5316 7760 5322 7812
rect 6546 7800 6552 7812
rect 6507 7772 6552 7800
rect 6546 7760 6552 7772
rect 6604 7760 6610 7812
rect 7006 7760 7012 7812
rect 7064 7760 7070 7812
rect 2685 7735 2743 7741
rect 2685 7701 2697 7735
rect 2731 7732 2743 7735
rect 5442 7732 5448 7744
rect 2731 7704 5448 7732
rect 2731 7701 2743 7704
rect 2685 7695 2743 7701
rect 5442 7692 5448 7704
rect 5500 7692 5506 7744
rect 10410 7732 10416 7744
rect 10371 7704 10416 7732
rect 10410 7692 10416 7704
rect 10468 7692 10474 7744
rect 1104 7642 11224 7664
rect 1104 7590 4323 7642
rect 4375 7590 4387 7642
rect 4439 7590 4451 7642
rect 4503 7590 4515 7642
rect 4567 7590 4579 7642
rect 4631 7590 7696 7642
rect 7748 7590 7760 7642
rect 7812 7590 7824 7642
rect 7876 7590 7888 7642
rect 7940 7590 7952 7642
rect 8004 7590 11224 7642
rect 1104 7568 11224 7590
rect 3050 7528 3056 7540
rect 2792 7500 3056 7528
rect 2792 7460 2820 7500
rect 3050 7488 3056 7500
rect 3108 7528 3114 7540
rect 3970 7528 3976 7540
rect 3108 7500 3976 7528
rect 3108 7488 3114 7500
rect 3970 7488 3976 7500
rect 4028 7488 4034 7540
rect 4890 7528 4896 7540
rect 4851 7500 4896 7528
rect 4890 7488 4896 7500
rect 4948 7488 4954 7540
rect 7929 7531 7987 7537
rect 7929 7497 7941 7531
rect 7975 7528 7987 7531
rect 8018 7528 8024 7540
rect 7975 7500 8024 7528
rect 7975 7497 7987 7500
rect 7929 7491 7987 7497
rect 8018 7488 8024 7500
rect 8076 7488 8082 7540
rect 2438 7432 2820 7460
rect 2869 7463 2927 7469
rect 2869 7429 2881 7463
rect 2915 7460 2927 7463
rect 4246 7460 4252 7472
rect 2915 7432 4252 7460
rect 2915 7429 2927 7432
rect 2869 7423 2927 7429
rect 4246 7420 4252 7432
rect 4304 7420 4310 7472
rect 4433 7463 4491 7469
rect 4433 7429 4445 7463
rect 4479 7460 4491 7463
rect 5074 7460 5080 7472
rect 4479 7432 5080 7460
rect 4479 7429 4491 7432
rect 4433 7423 4491 7429
rect 5074 7420 5080 7432
rect 5132 7460 5138 7472
rect 5132 7432 7696 7460
rect 5132 7420 5138 7432
rect 3142 7352 3148 7404
rect 3200 7392 3206 7404
rect 4525 7395 4583 7401
rect 3200 7364 3245 7392
rect 3200 7352 3206 7364
rect 4525 7361 4537 7395
rect 4571 7392 4583 7395
rect 7558 7392 7564 7404
rect 4571 7364 7564 7392
rect 4571 7361 4583 7364
rect 4525 7355 4583 7361
rect 7558 7352 7564 7364
rect 7616 7352 7622 7404
rect 4246 7324 4252 7336
rect 4207 7296 4252 7324
rect 4246 7284 4252 7296
rect 4304 7284 4310 7336
rect 7374 7324 7380 7336
rect 7335 7296 7380 7324
rect 7374 7284 7380 7296
rect 7432 7284 7438 7336
rect 7469 7327 7527 7333
rect 7469 7293 7481 7327
rect 7515 7324 7527 7327
rect 7668 7324 7696 7432
rect 8202 7420 8208 7472
rect 8260 7460 8266 7472
rect 8260 7432 9062 7460
rect 8260 7420 8266 7432
rect 8938 7324 8944 7336
rect 7515 7296 8944 7324
rect 7515 7293 7527 7296
rect 7469 7287 7527 7293
rect 8938 7284 8944 7296
rect 8996 7284 9002 7336
rect 10226 7324 10232 7336
rect 10187 7296 10232 7324
rect 10226 7284 10232 7296
rect 10284 7284 10290 7336
rect 10502 7324 10508 7336
rect 10463 7296 10508 7324
rect 10502 7284 10508 7296
rect 10560 7284 10566 7336
rect 5258 7216 5264 7268
rect 5316 7256 5322 7268
rect 8757 7259 8815 7265
rect 8757 7256 8769 7259
rect 5316 7228 8769 7256
rect 5316 7216 5322 7228
rect 8757 7225 8769 7228
rect 8803 7225 8815 7259
rect 8757 7219 8815 7225
rect 1394 7188 1400 7200
rect 1355 7160 1400 7188
rect 1394 7148 1400 7160
rect 1452 7148 1458 7200
rect 1104 7098 11224 7120
rect 1104 7046 2636 7098
rect 2688 7046 2700 7098
rect 2752 7046 2764 7098
rect 2816 7046 2828 7098
rect 2880 7046 2892 7098
rect 2944 7046 6010 7098
rect 6062 7046 6074 7098
rect 6126 7046 6138 7098
rect 6190 7046 6202 7098
rect 6254 7046 6266 7098
rect 6318 7046 9383 7098
rect 9435 7046 9447 7098
rect 9499 7046 9511 7098
rect 9563 7046 9575 7098
rect 9627 7046 9639 7098
rect 9691 7046 11224 7098
rect 1104 7024 11224 7046
rect 1486 6916 1492 6928
rect 1447 6888 1492 6916
rect 1486 6876 1492 6888
rect 1544 6876 1550 6928
rect 7006 6876 7012 6928
rect 7064 6916 7070 6928
rect 8202 6916 8208 6928
rect 7064 6888 8208 6916
rect 7064 6876 7070 6888
rect 8202 6876 8208 6888
rect 8260 6876 8266 6928
rect 6546 6808 6552 6860
rect 6604 6848 6610 6860
rect 7285 6851 7343 6857
rect 7285 6848 7297 6851
rect 6604 6820 7297 6848
rect 6604 6808 6610 6820
rect 7285 6817 7297 6820
rect 7331 6817 7343 6851
rect 7285 6811 7343 6817
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 2406 6780 2412 6792
rect 1719 6752 2412 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 2406 6740 2412 6752
rect 2464 6740 2470 6792
rect 3142 6740 3148 6792
rect 3200 6780 3206 6792
rect 5534 6780 5540 6792
rect 3200 6752 5540 6780
rect 3200 6740 3206 6752
rect 5534 6740 5540 6752
rect 5592 6740 5598 6792
rect 8110 6740 8116 6792
rect 8168 6780 8174 6792
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 8168 6752 9137 6780
rect 8168 6740 8174 6752
rect 9125 6749 9137 6752
rect 9171 6749 9183 6783
rect 9125 6743 9183 6749
rect 9309 6783 9367 6789
rect 9309 6749 9321 6783
rect 9355 6749 9367 6783
rect 9309 6743 9367 6749
rect 5810 6712 5816 6724
rect 5771 6684 5816 6712
rect 5810 6672 5816 6684
rect 5868 6672 5874 6724
rect 9324 6712 9352 6743
rect 9398 6740 9404 6792
rect 9456 6780 9462 6792
rect 9585 6783 9643 6789
rect 9585 6780 9597 6783
rect 9456 6752 9597 6780
rect 9456 6740 9462 6752
rect 9585 6749 9597 6752
rect 9631 6749 9643 6783
rect 9585 6743 9643 6749
rect 10134 6712 10140 6724
rect 6196 6684 6302 6712
rect 9324 6684 10140 6712
rect 2958 6604 2964 6656
rect 3016 6644 3022 6656
rect 3142 6644 3148 6656
rect 3016 6616 3148 6644
rect 3016 6604 3022 6616
rect 3142 6604 3148 6616
rect 3200 6604 3206 6656
rect 4062 6604 4068 6656
rect 4120 6644 4126 6656
rect 6196 6644 6224 6684
rect 10134 6672 10140 6684
rect 10192 6672 10198 6724
rect 4120 6616 6224 6644
rect 9769 6647 9827 6653
rect 4120 6604 4126 6616
rect 9769 6613 9781 6647
rect 9815 6644 9827 6647
rect 9858 6644 9864 6656
rect 9815 6616 9864 6644
rect 9815 6613 9827 6616
rect 9769 6607 9827 6613
rect 9858 6604 9864 6616
rect 9916 6604 9922 6656
rect 1104 6554 11224 6576
rect 1104 6502 4323 6554
rect 4375 6502 4387 6554
rect 4439 6502 4451 6554
rect 4503 6502 4515 6554
rect 4567 6502 4579 6554
rect 4631 6502 7696 6554
rect 7748 6502 7760 6554
rect 7812 6502 7824 6554
rect 7876 6502 7888 6554
rect 7940 6502 7952 6554
rect 8004 6502 11224 6554
rect 1104 6480 11224 6502
rect 5810 6440 5816 6452
rect 5771 6412 5816 6440
rect 5810 6400 5816 6412
rect 5868 6400 5874 6452
rect 6825 6443 6883 6449
rect 6825 6409 6837 6443
rect 6871 6440 6883 6443
rect 7558 6440 7564 6452
rect 6871 6412 7564 6440
rect 6871 6409 6883 6412
rect 6825 6403 6883 6409
rect 7558 6400 7564 6412
rect 7616 6400 7622 6452
rect 10137 6443 10195 6449
rect 10137 6409 10149 6443
rect 10183 6440 10195 6443
rect 10226 6440 10232 6452
rect 10183 6412 10232 6440
rect 10183 6409 10195 6412
rect 10137 6403 10195 6409
rect 10226 6400 10232 6412
rect 10284 6400 10290 6452
rect 1394 6332 1400 6384
rect 1452 6372 1458 6384
rect 2041 6375 2099 6381
rect 2041 6372 2053 6375
rect 1452 6344 2053 6372
rect 1452 6332 1458 6344
rect 2041 6341 2053 6344
rect 2087 6341 2099 6375
rect 2041 6335 2099 6341
rect 3050 6332 3056 6384
rect 3108 6332 3114 6384
rect 4062 6332 4068 6384
rect 4120 6372 4126 6384
rect 4120 6344 4830 6372
rect 4120 6332 4126 6344
rect 8202 6332 8208 6384
rect 8260 6372 8266 6384
rect 8260 6344 9154 6372
rect 8260 6332 8266 6344
rect 6917 6307 6975 6313
rect 6917 6273 6929 6307
rect 6963 6304 6975 6307
rect 7098 6304 7104 6316
rect 6963 6276 7104 6304
rect 6963 6273 6975 6276
rect 6917 6267 6975 6273
rect 7098 6264 7104 6276
rect 7156 6264 7162 6316
rect 1765 6239 1823 6245
rect 1765 6205 1777 6239
rect 1811 6236 1823 6239
rect 2774 6236 2780 6248
rect 1811 6208 2780 6236
rect 1811 6205 1823 6208
rect 1765 6199 1823 6205
rect 2774 6196 2780 6208
rect 2832 6236 2838 6248
rect 4065 6239 4123 6245
rect 4065 6236 4077 6239
rect 2832 6208 4077 6236
rect 2832 6196 2838 6208
rect 4065 6205 4077 6208
rect 4111 6205 4123 6239
rect 4338 6236 4344 6248
rect 4299 6208 4344 6236
rect 4065 6199 4123 6205
rect 4338 6196 4344 6208
rect 4396 6196 4402 6248
rect 8386 6236 8392 6248
rect 8347 6208 8392 6236
rect 8386 6196 8392 6208
rect 8444 6196 8450 6248
rect 8665 6239 8723 6245
rect 8665 6205 8677 6239
rect 8711 6236 8723 6239
rect 9030 6236 9036 6248
rect 8711 6208 9036 6236
rect 8711 6205 8723 6208
rect 8665 6199 8723 6205
rect 9030 6196 9036 6208
rect 9088 6236 9094 6248
rect 9398 6236 9404 6248
rect 9088 6208 9404 6236
rect 9088 6196 9094 6208
rect 9398 6196 9404 6208
rect 9456 6196 9462 6248
rect 3418 6060 3424 6112
rect 3476 6100 3482 6112
rect 3513 6103 3571 6109
rect 3513 6100 3525 6103
rect 3476 6072 3525 6100
rect 3476 6060 3482 6072
rect 3513 6069 3525 6072
rect 3559 6069 3571 6103
rect 3513 6063 3571 6069
rect 1104 6010 11224 6032
rect 1104 5958 2636 6010
rect 2688 5958 2700 6010
rect 2752 5958 2764 6010
rect 2816 5958 2828 6010
rect 2880 5958 2892 6010
rect 2944 5958 6010 6010
rect 6062 5958 6074 6010
rect 6126 5958 6138 6010
rect 6190 5958 6202 6010
rect 6254 5958 6266 6010
rect 6318 5958 9383 6010
rect 9435 5958 9447 6010
rect 9499 5958 9511 6010
rect 9563 5958 9575 6010
rect 9627 5958 9639 6010
rect 9691 5958 11224 6010
rect 1104 5936 11224 5958
rect 3789 5763 3847 5769
rect 3789 5760 3801 5763
rect 2700 5732 3801 5760
rect 2498 5692 2504 5704
rect 2459 5664 2504 5692
rect 2498 5652 2504 5664
rect 2556 5652 2562 5704
rect 2700 5701 2728 5732
rect 3789 5729 3801 5732
rect 3835 5729 3847 5763
rect 4154 5760 4160 5772
rect 3789 5723 3847 5729
rect 3988 5732 4160 5760
rect 2685 5695 2743 5701
rect 2685 5661 2697 5695
rect 2731 5661 2743 5695
rect 2685 5655 2743 5661
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5692 3019 5695
rect 3694 5692 3700 5704
rect 3007 5664 3700 5692
rect 3007 5661 3019 5664
rect 2961 5655 3019 5661
rect 3694 5652 3700 5664
rect 3752 5652 3758 5704
rect 3988 5701 4016 5732
rect 4154 5720 4160 5732
rect 4212 5760 4218 5772
rect 4338 5760 4344 5772
rect 4212 5732 4344 5760
rect 4212 5720 4218 5732
rect 4338 5720 4344 5732
rect 4396 5720 4402 5772
rect 6914 5720 6920 5772
rect 6972 5760 6978 5772
rect 8110 5760 8116 5772
rect 6972 5732 8116 5760
rect 6972 5720 6978 5732
rect 8110 5720 8116 5732
rect 8168 5720 8174 5772
rect 9030 5760 9036 5772
rect 8991 5732 9036 5760
rect 9030 5720 9036 5732
rect 9088 5720 9094 5772
rect 3973 5695 4031 5701
rect 3973 5661 3985 5695
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 4249 5695 4307 5701
rect 4249 5661 4261 5695
rect 4295 5661 4307 5695
rect 4249 5655 4307 5661
rect 4433 5695 4491 5701
rect 4433 5661 4445 5695
rect 4479 5692 4491 5695
rect 4798 5692 4804 5704
rect 4479 5664 4804 5692
rect 4479 5661 4491 5664
rect 4433 5655 4491 5661
rect 3418 5584 3424 5636
rect 3476 5624 3482 5636
rect 4264 5624 4292 5655
rect 4798 5652 4804 5664
rect 4856 5652 4862 5704
rect 7006 5652 7012 5704
rect 7064 5652 7070 5704
rect 8386 5652 8392 5704
rect 8444 5692 8450 5704
rect 8444 5664 8489 5692
rect 8444 5652 8450 5664
rect 8938 5652 8944 5704
rect 8996 5692 9002 5704
rect 9217 5695 9275 5701
rect 9217 5692 9229 5695
rect 8996 5664 9229 5692
rect 8996 5652 9002 5664
rect 9217 5661 9229 5664
rect 9263 5661 9275 5695
rect 9217 5655 9275 5661
rect 3476 5596 4292 5624
rect 3476 5584 3482 5596
rect 3142 5556 3148 5568
rect 3103 5528 3148 5556
rect 3142 5516 3148 5528
rect 3200 5516 3206 5568
rect 6641 5559 6699 5565
rect 6641 5525 6653 5559
rect 6687 5556 6699 5559
rect 7098 5556 7104 5568
rect 6687 5528 7104 5556
rect 6687 5525 6699 5528
rect 6641 5519 6699 5525
rect 7098 5516 7104 5528
rect 7156 5556 7162 5568
rect 8110 5556 8116 5568
rect 7156 5528 8116 5556
rect 7156 5516 7162 5528
rect 8110 5516 8116 5528
rect 8168 5556 8174 5568
rect 9309 5559 9367 5565
rect 9309 5556 9321 5559
rect 8168 5528 9321 5556
rect 8168 5516 8174 5528
rect 9309 5525 9321 5528
rect 9355 5525 9367 5559
rect 9309 5519 9367 5525
rect 9677 5559 9735 5565
rect 9677 5525 9689 5559
rect 9723 5556 9735 5559
rect 9766 5556 9772 5568
rect 9723 5528 9772 5556
rect 9723 5525 9735 5528
rect 9677 5519 9735 5525
rect 9766 5516 9772 5528
rect 9824 5516 9830 5568
rect 1104 5466 11224 5488
rect 1104 5414 4323 5466
rect 4375 5414 4387 5466
rect 4439 5414 4451 5466
rect 4503 5414 4515 5466
rect 4567 5414 4579 5466
rect 4631 5414 7696 5466
rect 7748 5414 7760 5466
rect 7812 5414 7824 5466
rect 7876 5414 7888 5466
rect 7940 5414 7952 5466
rect 8004 5414 11224 5466
rect 1104 5392 11224 5414
rect 2314 5312 2320 5364
rect 2372 5352 2378 5364
rect 3050 5352 3056 5364
rect 2372 5324 3056 5352
rect 2372 5312 2378 5324
rect 3050 5312 3056 5324
rect 3108 5352 3114 5364
rect 4062 5352 4068 5364
rect 3108 5324 4068 5352
rect 3108 5312 3114 5324
rect 3145 5287 3203 5293
rect 3145 5253 3157 5287
rect 3191 5284 3203 5287
rect 3418 5284 3424 5296
rect 3191 5256 3424 5284
rect 3191 5253 3203 5256
rect 3145 5247 3203 5253
rect 3418 5244 3424 5256
rect 3476 5244 3482 5296
rect 3528 5284 3556 5324
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 4154 5312 4160 5364
rect 4212 5352 4218 5364
rect 4617 5355 4675 5361
rect 4617 5352 4629 5355
rect 4212 5324 4629 5352
rect 4212 5312 4218 5324
rect 4617 5321 4629 5324
rect 4663 5321 4675 5355
rect 7006 5352 7012 5364
rect 4617 5315 4675 5321
rect 6564 5324 7012 5352
rect 3528 5256 3634 5284
rect 5442 5244 5448 5296
rect 5500 5284 5506 5296
rect 6564 5284 6592 5324
rect 7006 5312 7012 5324
rect 7064 5352 7070 5364
rect 8757 5355 8815 5361
rect 7064 5324 8248 5352
rect 7064 5312 7070 5324
rect 8220 5296 8248 5324
rect 8757 5321 8769 5355
rect 8803 5352 8815 5355
rect 8938 5352 8944 5364
rect 8803 5324 8944 5352
rect 8803 5321 8815 5324
rect 8757 5315 8815 5321
rect 8938 5312 8944 5324
rect 8996 5312 9002 5364
rect 7837 5287 7895 5293
rect 5500 5256 6670 5284
rect 5500 5244 5506 5256
rect 7837 5253 7849 5287
rect 7883 5284 7895 5287
rect 8110 5284 8116 5296
rect 7883 5256 8116 5284
rect 7883 5253 7895 5256
rect 7837 5247 7895 5253
rect 8110 5244 8116 5256
rect 8168 5244 8174 5296
rect 8202 5244 8208 5296
rect 8260 5284 8266 5296
rect 8260 5256 9062 5284
rect 8260 5244 8266 5256
rect 10134 5244 10140 5296
rect 10192 5284 10198 5296
rect 10229 5287 10287 5293
rect 10229 5284 10241 5287
rect 10192 5256 10241 5284
rect 10192 5244 10198 5256
rect 10229 5253 10241 5256
rect 10275 5284 10287 5287
rect 10318 5284 10324 5296
rect 10275 5256 10324 5284
rect 10275 5253 10287 5256
rect 10229 5247 10287 5253
rect 10318 5244 10324 5256
rect 10376 5244 10382 5296
rect 2866 5216 2872 5228
rect 2827 5188 2872 5216
rect 2866 5176 2872 5188
rect 2924 5176 2930 5228
rect 5350 5216 5356 5228
rect 5311 5188 5356 5216
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 5626 5216 5632 5228
rect 5587 5188 5632 5216
rect 5626 5176 5632 5188
rect 5684 5176 5690 5228
rect 5718 5176 5724 5228
rect 5776 5216 5782 5228
rect 5813 5219 5871 5225
rect 5813 5216 5825 5219
rect 5776 5188 5825 5216
rect 5776 5176 5782 5188
rect 5813 5185 5825 5188
rect 5859 5185 5871 5219
rect 5813 5179 5871 5185
rect 10502 5176 10508 5228
rect 10560 5216 10566 5228
rect 10560 5188 10605 5216
rect 10560 5176 10566 5188
rect 6638 5108 6644 5160
rect 6696 5148 6702 5160
rect 8113 5151 8171 5157
rect 8113 5148 8125 5151
rect 6696 5120 8125 5148
rect 6696 5108 6702 5120
rect 8113 5117 8125 5120
rect 8159 5148 8171 5151
rect 8386 5148 8392 5160
rect 8159 5120 8392 5148
rect 8159 5117 8171 5120
rect 8113 5111 8171 5117
rect 8386 5108 8392 5120
rect 8444 5148 8450 5160
rect 10520 5148 10548 5176
rect 8444 5120 10548 5148
rect 8444 5108 8450 5120
rect 4798 4972 4804 5024
rect 4856 5012 4862 5024
rect 5169 5015 5227 5021
rect 5169 5012 5181 5015
rect 4856 4984 5181 5012
rect 4856 4972 4862 4984
rect 5169 4981 5181 4984
rect 5215 4981 5227 5015
rect 5169 4975 5227 4981
rect 6365 5015 6423 5021
rect 6365 4981 6377 5015
rect 6411 5012 6423 5015
rect 7190 5012 7196 5024
rect 6411 4984 7196 5012
rect 6411 4981 6423 4984
rect 6365 4975 6423 4981
rect 7190 4972 7196 4984
rect 7248 4972 7254 5024
rect 1104 4922 11224 4944
rect 1104 4870 2636 4922
rect 2688 4870 2700 4922
rect 2752 4870 2764 4922
rect 2816 4870 2828 4922
rect 2880 4870 2892 4922
rect 2944 4870 6010 4922
rect 6062 4870 6074 4922
rect 6126 4870 6138 4922
rect 6190 4870 6202 4922
rect 6254 4870 6266 4922
rect 6318 4870 9383 4922
rect 9435 4870 9447 4922
rect 9499 4870 9511 4922
rect 9563 4870 9575 4922
rect 9627 4870 9639 4922
rect 9691 4870 11224 4922
rect 1104 4848 11224 4870
rect 1397 4811 1455 4817
rect 1397 4777 1409 4811
rect 1443 4808 1455 4811
rect 2498 4808 2504 4820
rect 1443 4780 2504 4808
rect 1443 4777 1455 4780
rect 1397 4771 1455 4777
rect 2498 4768 2504 4780
rect 2556 4768 2562 4820
rect 3694 4768 3700 4820
rect 3752 4808 3758 4820
rect 3789 4811 3847 4817
rect 3789 4808 3801 4811
rect 3752 4780 3801 4808
rect 3752 4768 3758 4780
rect 3789 4777 3801 4780
rect 3835 4777 3847 4811
rect 3789 4771 3847 4777
rect 5626 4768 5632 4820
rect 5684 4808 5690 4820
rect 6181 4811 6239 4817
rect 6181 4808 6193 4811
rect 5684 4780 6193 4808
rect 5684 4768 5690 4780
rect 6181 4777 6193 4780
rect 6227 4777 6239 4811
rect 6181 4771 6239 4777
rect 3142 4700 3148 4752
rect 3200 4700 3206 4752
rect 4890 4700 4896 4752
rect 4948 4740 4954 4752
rect 4948 4712 6914 4740
rect 4948 4700 4954 4712
rect 2869 4675 2927 4681
rect 2869 4641 2881 4675
rect 2915 4672 2927 4675
rect 3160 4672 3188 4700
rect 2915 4644 3188 4672
rect 2915 4641 2927 4644
rect 2869 4635 2927 4641
rect 4154 4632 4160 4684
rect 4212 4672 4218 4684
rect 4341 4675 4399 4681
rect 4341 4672 4353 4675
rect 4212 4644 4353 4672
rect 4212 4632 4218 4644
rect 4341 4641 4353 4644
rect 4387 4641 4399 4675
rect 4341 4635 4399 4641
rect 5166 4632 5172 4684
rect 5224 4672 5230 4684
rect 5537 4675 5595 4681
rect 5537 4672 5549 4675
rect 5224 4644 5549 4672
rect 5224 4632 5230 4644
rect 5537 4641 5549 4644
rect 5583 4641 5595 4675
rect 6886 4672 6914 4712
rect 5537 4635 5595 4641
rect 6840 4644 8064 4672
rect 3145 4607 3203 4613
rect 3145 4573 3157 4607
rect 3191 4573 3203 4607
rect 3145 4567 3203 4573
rect 5445 4607 5503 4613
rect 5445 4573 5457 4607
rect 5491 4604 5503 4607
rect 5718 4604 5724 4616
rect 5491 4576 5724 4604
rect 5491 4573 5503 4576
rect 5445 4567 5503 4573
rect 2314 4496 2320 4548
rect 2372 4496 2378 4548
rect 2958 4496 2964 4548
rect 3016 4536 3022 4548
rect 3160 4536 3188 4567
rect 5718 4564 5724 4576
rect 5776 4564 5782 4616
rect 6362 4604 6368 4616
rect 6323 4576 6368 4604
rect 6362 4564 6368 4576
rect 6420 4564 6426 4616
rect 6840 4613 6868 4644
rect 6641 4607 6699 4613
rect 6641 4573 6653 4607
rect 6687 4573 6699 4607
rect 6641 4567 6699 4573
rect 6825 4607 6883 4613
rect 6825 4573 6837 4607
rect 6871 4573 6883 4607
rect 6825 4567 6883 4573
rect 3016 4508 3188 4536
rect 4157 4539 4215 4545
rect 3016 4496 3022 4508
rect 4157 4505 4169 4539
rect 4203 4536 4215 4539
rect 5534 4536 5540 4548
rect 4203 4508 5540 4536
rect 4203 4505 4215 4508
rect 4157 4499 4215 4505
rect 5534 4496 5540 4508
rect 5592 4496 5598 4548
rect 6656 4536 6684 4567
rect 7466 4564 7472 4616
rect 7524 4604 7530 4616
rect 8036 4613 8064 4644
rect 8202 4632 8208 4684
rect 8260 4672 8266 4684
rect 9306 4672 9312 4684
rect 8260 4644 9312 4672
rect 8260 4632 8266 4644
rect 9306 4632 9312 4644
rect 9364 4632 9370 4684
rect 7561 4607 7619 4613
rect 7561 4604 7573 4607
rect 7524 4576 7573 4604
rect 7524 4564 7530 4576
rect 7561 4573 7573 4576
rect 7607 4573 7619 4607
rect 7561 4567 7619 4573
rect 7837 4607 7895 4613
rect 7837 4573 7849 4607
rect 7883 4573 7895 4607
rect 7837 4567 7895 4573
rect 8021 4607 8079 4613
rect 8021 4573 8033 4607
rect 8067 4573 8079 4607
rect 10502 4604 10508 4616
rect 10463 4576 10508 4604
rect 8021 4567 8079 4573
rect 7190 4536 7196 4548
rect 6656 4508 7196 4536
rect 7190 4496 7196 4508
rect 7248 4496 7254 4548
rect 7852 4536 7880 4567
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 8202 4536 8208 4548
rect 7852 4508 8208 4536
rect 8202 4496 8208 4508
rect 8260 4496 8266 4548
rect 4246 4468 4252 4480
rect 4207 4440 4252 4468
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 4982 4468 4988 4480
rect 4943 4440 4988 4468
rect 4982 4428 4988 4440
rect 5040 4428 5046 4480
rect 5258 4428 5264 4480
rect 5316 4468 5322 4480
rect 5353 4471 5411 4477
rect 5353 4468 5365 4471
rect 5316 4440 5365 4468
rect 5316 4428 5322 4440
rect 5353 4437 5365 4440
rect 5399 4437 5411 4471
rect 5353 4431 5411 4437
rect 6914 4428 6920 4480
rect 6972 4468 6978 4480
rect 7377 4471 7435 4477
rect 7377 4468 7389 4471
rect 6972 4440 7389 4468
rect 6972 4428 6978 4440
rect 7377 4437 7389 4440
rect 7423 4437 7435 4471
rect 7377 4431 7435 4437
rect 1104 4378 11224 4400
rect 1104 4326 4323 4378
rect 4375 4326 4387 4378
rect 4439 4326 4451 4378
rect 4503 4326 4515 4378
rect 4567 4326 4579 4378
rect 4631 4326 7696 4378
rect 7748 4326 7760 4378
rect 7812 4326 7824 4378
rect 7876 4326 7888 4378
rect 7940 4326 7952 4378
rect 8004 4326 11224 4378
rect 1104 4304 11224 4326
rect 5077 4267 5135 4273
rect 5077 4233 5089 4267
rect 5123 4264 5135 4267
rect 5350 4264 5356 4276
rect 5123 4236 5356 4264
rect 5123 4233 5135 4236
rect 5077 4227 5135 4233
rect 5350 4224 5356 4236
rect 5408 4224 5414 4276
rect 5445 4267 5503 4273
rect 5445 4233 5457 4267
rect 5491 4264 5503 4267
rect 5534 4264 5540 4276
rect 5491 4236 5540 4264
rect 5491 4233 5503 4236
rect 5445 4227 5503 4233
rect 5534 4224 5540 4236
rect 5592 4264 5598 4276
rect 7466 4264 7472 4276
rect 5592 4236 7472 4264
rect 5592 4224 5598 4236
rect 7466 4224 7472 4236
rect 7524 4224 7530 4276
rect 10318 4224 10324 4276
rect 10376 4264 10382 4276
rect 10505 4267 10563 4273
rect 10505 4264 10517 4267
rect 10376 4236 10517 4264
rect 10376 4224 10382 4236
rect 10505 4233 10517 4236
rect 10551 4233 10563 4267
rect 10505 4227 10563 4233
rect 4154 4156 4160 4208
rect 4212 4196 4218 4208
rect 4212 4168 6670 4196
rect 4212 4156 4218 4168
rect 5460 4140 5488 4168
rect 9306 4156 9312 4208
rect 9364 4196 9370 4208
rect 9364 4168 9522 4196
rect 9364 4156 9370 4168
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4097 1731 4131
rect 2130 4128 2136 4140
rect 2091 4100 2136 4128
rect 1673 4091 1731 4097
rect 1688 4060 1716 4091
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4128 4307 4131
rect 4982 4128 4988 4140
rect 4295 4100 4988 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 5442 4088 5448 4140
rect 5500 4088 5506 4140
rect 2222 4060 2228 4072
rect 1688 4032 2228 4060
rect 2222 4020 2228 4032
rect 2280 4020 2286 4072
rect 4338 4020 4344 4072
rect 4396 4060 4402 4072
rect 5074 4060 5080 4072
rect 4396 4032 5080 4060
rect 4396 4020 4402 4032
rect 5074 4020 5080 4032
rect 5132 4060 5138 4072
rect 5537 4063 5595 4069
rect 5537 4060 5549 4063
rect 5132 4032 5549 4060
rect 5132 4020 5138 4032
rect 5537 4029 5549 4032
rect 5583 4029 5595 4063
rect 5537 4023 5595 4029
rect 5721 4063 5779 4069
rect 5721 4029 5733 4063
rect 5767 4060 5779 4063
rect 6362 4060 6368 4072
rect 5767 4032 6368 4060
rect 5767 4029 5779 4032
rect 5721 4023 5779 4029
rect 6362 4020 6368 4032
rect 6420 4020 6426 4072
rect 7190 4020 7196 4072
rect 7248 4060 7254 4072
rect 7837 4063 7895 4069
rect 7837 4060 7849 4063
rect 7248 4032 7849 4060
rect 7248 4020 7254 4032
rect 7837 4029 7849 4032
rect 7883 4029 7895 4063
rect 8113 4063 8171 4069
rect 8113 4060 8125 4063
rect 7837 4023 7895 4029
rect 8036 4032 8125 4060
rect 2038 3952 2044 4004
rect 2096 3992 2102 4004
rect 5166 3992 5172 4004
rect 2096 3964 5172 3992
rect 2096 3952 2102 3964
rect 5166 3952 5172 3964
rect 5224 3952 5230 4004
rect 1486 3924 1492 3936
rect 1447 3896 1492 3924
rect 1486 3884 1492 3896
rect 1544 3884 1550 3936
rect 2317 3927 2375 3933
rect 2317 3893 2329 3927
rect 2363 3924 2375 3927
rect 2498 3924 2504 3936
rect 2363 3896 2504 3924
rect 2363 3893 2375 3896
rect 2317 3887 2375 3893
rect 2498 3884 2504 3896
rect 2556 3884 2562 3936
rect 3878 3884 3884 3936
rect 3936 3924 3942 3936
rect 4065 3927 4123 3933
rect 4065 3924 4077 3927
rect 3936 3896 4077 3924
rect 3936 3884 3942 3896
rect 4065 3893 4077 3896
rect 4111 3893 4123 3927
rect 6362 3924 6368 3936
rect 6323 3896 6368 3924
rect 4065 3887 4123 3893
rect 6362 3884 6368 3896
rect 6420 3884 6426 3936
rect 6638 3884 6644 3936
rect 6696 3924 6702 3936
rect 8036 3924 8064 4032
rect 8113 4029 8125 4032
rect 8159 4060 8171 4063
rect 8757 4063 8815 4069
rect 8757 4060 8769 4063
rect 8159 4032 8769 4060
rect 8159 4029 8171 4032
rect 8113 4023 8171 4029
rect 8757 4029 8769 4032
rect 8803 4029 8815 4063
rect 9030 4060 9036 4072
rect 8991 4032 9036 4060
rect 8757 4023 8815 4029
rect 9030 4020 9036 4032
rect 9088 4020 9094 4072
rect 6696 3896 8064 3924
rect 6696 3884 6702 3896
rect 1104 3834 11224 3856
rect 1104 3782 2636 3834
rect 2688 3782 2700 3834
rect 2752 3782 2764 3834
rect 2816 3782 2828 3834
rect 2880 3782 2892 3834
rect 2944 3782 6010 3834
rect 6062 3782 6074 3834
rect 6126 3782 6138 3834
rect 6190 3782 6202 3834
rect 6254 3782 6266 3834
rect 6318 3782 9383 3834
rect 9435 3782 9447 3834
rect 9499 3782 9511 3834
rect 9563 3782 9575 3834
rect 9627 3782 9639 3834
rect 9691 3782 11224 3834
rect 1104 3760 11224 3782
rect 2130 3680 2136 3732
rect 2188 3720 2194 3732
rect 2593 3723 2651 3729
rect 2593 3720 2605 3723
rect 2188 3692 2605 3720
rect 2188 3680 2194 3692
rect 2593 3689 2605 3692
rect 2639 3689 2651 3723
rect 2593 3683 2651 3689
rect 5718 3680 5724 3732
rect 5776 3720 5782 3732
rect 5813 3723 5871 3729
rect 5813 3720 5825 3723
rect 5776 3692 5825 3720
rect 5776 3680 5782 3692
rect 5813 3689 5825 3692
rect 5859 3689 5871 3723
rect 5813 3683 5871 3689
rect 9766 3652 9772 3664
rect 9324 3624 9772 3652
rect 2038 3584 2044 3596
rect 1999 3556 2044 3584
rect 2038 3544 2044 3556
rect 2096 3544 2102 3596
rect 2133 3587 2191 3593
rect 2133 3553 2145 3587
rect 2179 3584 2191 3587
rect 2406 3584 2412 3596
rect 2179 3556 2412 3584
rect 2179 3553 2191 3556
rect 2133 3547 2191 3553
rect 2406 3544 2412 3556
rect 2464 3544 2470 3596
rect 2958 3544 2964 3596
rect 3016 3584 3022 3596
rect 4062 3584 4068 3596
rect 3016 3556 4068 3584
rect 3016 3544 3022 3556
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 4341 3587 4399 3593
rect 4341 3553 4353 3587
rect 4387 3584 4399 3587
rect 4798 3584 4804 3596
rect 4387 3556 4804 3584
rect 4387 3553 4399 3556
rect 4341 3547 4399 3553
rect 4798 3544 4804 3556
rect 4856 3544 4862 3596
rect 6917 3587 6975 3593
rect 6917 3553 6929 3587
rect 6963 3584 6975 3587
rect 9125 3587 9183 3593
rect 9125 3584 9137 3587
rect 6963 3556 9137 3584
rect 6963 3553 6975 3556
rect 6917 3547 6975 3553
rect 9125 3553 9137 3556
rect 9171 3553 9183 3587
rect 9125 3547 9183 3553
rect 6638 3516 6644 3528
rect 6599 3488 6644 3516
rect 6638 3476 6644 3488
rect 6696 3476 6702 3528
rect 8018 3476 8024 3528
rect 8076 3476 8082 3528
rect 9324 3525 9352 3624
rect 9766 3612 9772 3624
rect 9824 3612 9830 3664
rect 9858 3584 9864 3596
rect 9600 3556 9864 3584
rect 9600 3525 9628 3556
rect 9858 3544 9864 3556
rect 9916 3544 9922 3596
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3485 9367 3519
rect 9309 3479 9367 3485
rect 9585 3519 9643 3525
rect 9585 3485 9597 3519
rect 9631 3485 9643 3519
rect 9585 3479 9643 3485
rect 9769 3519 9827 3525
rect 9769 3485 9781 3519
rect 9815 3516 9827 3519
rect 9950 3516 9956 3528
rect 9815 3488 9956 3516
rect 9815 3485 9827 3488
rect 9769 3479 9827 3485
rect 4172 3420 4830 3448
rect 4172 3392 4200 3420
rect 2222 3340 2228 3392
rect 2280 3380 2286 3392
rect 2280 3352 2325 3380
rect 2280 3340 2286 3352
rect 4154 3340 4160 3392
rect 4212 3340 4218 3392
rect 8389 3383 8447 3389
rect 8389 3349 8401 3383
rect 8435 3380 8447 3383
rect 9784 3380 9812 3479
rect 9950 3476 9956 3488
rect 10008 3476 10014 3528
rect 8435 3352 9812 3380
rect 8435 3349 8447 3352
rect 8389 3343 8447 3349
rect 1104 3290 11224 3312
rect 1104 3238 4323 3290
rect 4375 3238 4387 3290
rect 4439 3238 4451 3290
rect 4503 3238 4515 3290
rect 4567 3238 4579 3290
rect 4631 3238 7696 3290
rect 7748 3238 7760 3290
rect 7812 3238 7824 3290
rect 7876 3238 7888 3290
rect 7940 3238 7952 3290
rect 8004 3238 11224 3290
rect 1104 3216 11224 3238
rect 1397 3179 1455 3185
rect 1397 3145 1409 3179
rect 1443 3176 1455 3179
rect 2222 3176 2228 3188
rect 1443 3148 2228 3176
rect 1443 3145 1455 3148
rect 1397 3139 1455 3145
rect 2222 3136 2228 3148
rect 2280 3136 2286 3188
rect 2498 3136 2504 3188
rect 2556 3136 2562 3188
rect 5258 3136 5264 3188
rect 5316 3176 5322 3188
rect 5353 3179 5411 3185
rect 5353 3176 5365 3179
rect 5316 3148 5365 3176
rect 5316 3136 5322 3148
rect 5353 3145 5365 3148
rect 5399 3145 5411 3179
rect 5353 3139 5411 3145
rect 8941 3179 8999 3185
rect 8941 3145 8953 3179
rect 8987 3176 8999 3179
rect 9030 3176 9036 3188
rect 8987 3148 9036 3176
rect 8987 3145 8999 3148
rect 8941 3139 8999 3145
rect 2314 3068 2320 3120
rect 2372 3068 2378 3120
rect 2516 3108 2544 3136
rect 2869 3111 2927 3117
rect 2869 3108 2881 3111
rect 2516 3080 2881 3108
rect 2869 3077 2881 3080
rect 2915 3077 2927 3111
rect 2869 3071 2927 3077
rect 2958 3068 2964 3120
rect 3016 3108 3022 3120
rect 3878 3108 3884 3120
rect 3016 3080 3188 3108
rect 3839 3080 3884 3108
rect 3016 3068 3022 3080
rect 3160 3049 3188 3080
rect 3878 3068 3884 3080
rect 3936 3068 3942 3120
rect 4154 3068 4160 3120
rect 4212 3108 4218 3120
rect 4212 3080 4370 3108
rect 4212 3068 4218 3080
rect 3145 3043 3203 3049
rect 3145 3009 3157 3043
rect 3191 3040 3203 3043
rect 3605 3043 3663 3049
rect 3605 3040 3617 3043
rect 3191 3012 3617 3040
rect 3191 3009 3203 3012
rect 3145 3003 3203 3009
rect 3605 3009 3617 3012
rect 3651 3009 3663 3043
rect 5368 3040 5396 3139
rect 9030 3136 9036 3148
rect 9088 3136 9094 3188
rect 6362 3068 6368 3120
rect 6420 3108 6426 3120
rect 7469 3111 7527 3117
rect 7469 3108 7481 3111
rect 6420 3080 7481 3108
rect 6420 3068 6426 3080
rect 7469 3077 7481 3080
rect 7515 3077 7527 3111
rect 7469 3071 7527 3077
rect 8018 3068 8024 3120
rect 8076 3068 8082 3120
rect 6457 3043 6515 3049
rect 6457 3040 6469 3043
rect 5368 3012 6469 3040
rect 3605 3003 3663 3009
rect 6457 3009 6469 3012
rect 6503 3009 6515 3043
rect 6457 3003 6515 3009
rect 6638 3000 6644 3052
rect 6696 3040 6702 3052
rect 7193 3043 7251 3049
rect 7193 3040 7205 3043
rect 6696 3012 7205 3040
rect 6696 3000 6702 3012
rect 7193 3009 7205 3012
rect 7239 3009 7251 3043
rect 7193 3003 7251 3009
rect 6454 2796 6460 2848
rect 6512 2836 6518 2848
rect 6641 2839 6699 2845
rect 6641 2836 6653 2839
rect 6512 2808 6653 2836
rect 6512 2796 6518 2808
rect 6641 2805 6653 2808
rect 6687 2805 6699 2839
rect 6641 2799 6699 2805
rect 1104 2746 11224 2768
rect 1104 2694 2636 2746
rect 2688 2694 2700 2746
rect 2752 2694 2764 2746
rect 2816 2694 2828 2746
rect 2880 2694 2892 2746
rect 2944 2694 6010 2746
rect 6062 2694 6074 2746
rect 6126 2694 6138 2746
rect 6190 2694 6202 2746
rect 6254 2694 6266 2746
rect 6318 2694 9383 2746
rect 9435 2694 9447 2746
rect 9499 2694 9511 2746
rect 9563 2694 9575 2746
rect 9627 2694 9639 2746
rect 9691 2694 11224 2746
rect 1104 2672 11224 2694
rect 8202 2592 8208 2644
rect 8260 2632 8266 2644
rect 8389 2635 8447 2641
rect 8389 2632 8401 2635
rect 8260 2604 8401 2632
rect 8260 2592 8266 2604
rect 8389 2601 8401 2604
rect 8435 2601 8447 2635
rect 8389 2595 8447 2601
rect 2041 2567 2099 2573
rect 2041 2533 2053 2567
rect 2087 2564 2099 2567
rect 4246 2564 4252 2576
rect 2087 2536 4252 2564
rect 2087 2533 2099 2536
rect 2041 2527 2099 2533
rect 4246 2524 4252 2536
rect 4304 2524 4310 2576
rect 4154 2496 4160 2508
rect 4115 2468 4160 2496
rect 4154 2456 4160 2468
rect 4212 2496 4218 2508
rect 6638 2496 6644 2508
rect 4212 2468 6644 2496
rect 4212 2456 4218 2468
rect 6638 2456 6644 2468
rect 6696 2456 6702 2508
rect 6914 2456 6920 2508
rect 6972 2496 6978 2508
rect 6972 2468 7017 2496
rect 6972 2456 6978 2468
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 3292 2400 3801 2428
rect 3292 2388 3298 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 8018 2388 8024 2440
rect 8076 2388 8082 2440
rect 8404 2428 8432 2595
rect 9493 2431 9551 2437
rect 9493 2428 9505 2431
rect 8404 2400 9505 2428
rect 9493 2397 9505 2400
rect 9539 2397 9551 2431
rect 9493 2391 9551 2397
rect 9950 2388 9956 2440
rect 10008 2428 10014 2440
rect 10229 2431 10287 2437
rect 10229 2428 10241 2431
rect 10008 2400 10241 2428
rect 10008 2388 10014 2400
rect 10229 2397 10241 2400
rect 10275 2397 10287 2431
rect 10229 2391 10287 2397
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1857 2363 1915 2369
rect 1857 2360 1869 2363
rect 72 2332 1869 2360
rect 72 2320 78 2332
rect 1857 2329 1869 2332
rect 1903 2329 1915 2363
rect 1857 2323 1915 2329
rect 9674 2292 9680 2304
rect 9635 2264 9680 2292
rect 9674 2252 9680 2264
rect 9732 2252 9738 2304
rect 10410 2292 10416 2304
rect 10371 2264 10416 2292
rect 10410 2252 10416 2264
rect 10468 2252 10474 2304
rect 1104 2202 11224 2224
rect 1104 2150 4323 2202
rect 4375 2150 4387 2202
rect 4439 2150 4451 2202
rect 4503 2150 4515 2202
rect 4567 2150 4579 2202
rect 4631 2150 7696 2202
rect 7748 2150 7760 2202
rect 7812 2150 7824 2202
rect 7876 2150 7888 2202
rect 7940 2150 7952 2202
rect 8004 2150 11224 2202
rect 1104 2128 11224 2150
<< via1 >>
rect 4323 11942 4375 11994
rect 4387 11942 4439 11994
rect 4451 11942 4503 11994
rect 4515 11942 4567 11994
rect 4579 11942 4631 11994
rect 7696 11942 7748 11994
rect 7760 11942 7812 11994
rect 7824 11942 7876 11994
rect 7888 11942 7940 11994
rect 7952 11942 8004 11994
rect 1492 11883 1544 11892
rect 1492 11849 1501 11883
rect 1501 11849 1535 11883
rect 1535 11849 1544 11883
rect 1492 11840 1544 11849
rect 5816 11840 5868 11892
rect 9220 11883 9272 11892
rect 9220 11849 9229 11883
rect 9229 11849 9263 11883
rect 9263 11849 9272 11883
rect 9220 11840 9272 11849
rect 12256 11840 12308 11892
rect 2504 11704 2556 11756
rect 2688 11747 2740 11756
rect 2688 11713 2697 11747
rect 2697 11713 2731 11747
rect 2731 11713 2740 11747
rect 2688 11704 2740 11713
rect 5724 11704 5776 11756
rect 8944 11704 8996 11756
rect 9036 11704 9088 11756
rect 10140 11704 10192 11756
rect 3700 11568 3752 11620
rect 2964 11500 3016 11552
rect 6552 11500 6604 11552
rect 7564 11500 7616 11552
rect 2636 11398 2688 11450
rect 2700 11398 2752 11450
rect 2764 11398 2816 11450
rect 2828 11398 2880 11450
rect 2892 11398 2944 11450
rect 6010 11398 6062 11450
rect 6074 11398 6126 11450
rect 6138 11398 6190 11450
rect 6202 11398 6254 11450
rect 6266 11398 6318 11450
rect 9383 11398 9435 11450
rect 9447 11398 9499 11450
rect 9511 11398 9563 11450
rect 9575 11398 9627 11450
rect 9639 11398 9691 11450
rect 10416 11271 10468 11280
rect 10416 11237 10425 11271
rect 10425 11237 10459 11271
rect 10459 11237 10468 11271
rect 10416 11228 10468 11237
rect 1768 11135 1820 11144
rect 1768 11101 1777 11135
rect 1777 11101 1811 11135
rect 1811 11101 1820 11135
rect 1768 11092 1820 11101
rect 5908 11135 5960 11144
rect 5908 11101 5917 11135
rect 5917 11101 5951 11135
rect 5951 11101 5960 11135
rect 5908 11092 5960 11101
rect 10140 11160 10192 11212
rect 10048 11092 10100 11144
rect 10232 11135 10284 11144
rect 10232 11101 10241 11135
rect 10241 11101 10275 11135
rect 10275 11101 10284 11135
rect 10232 11092 10284 11101
rect 4068 11024 4120 11076
rect 5632 11067 5684 11076
rect 5632 11033 5641 11067
rect 5641 11033 5675 11067
rect 5675 11033 5684 11067
rect 5632 11024 5684 11033
rect 8668 11024 8720 11076
rect 4160 10999 4212 11008
rect 4160 10965 4169 10999
rect 4169 10965 4203 10999
rect 4203 10965 4212 10999
rect 4160 10956 4212 10965
rect 4323 10854 4375 10906
rect 4387 10854 4439 10906
rect 4451 10854 4503 10906
rect 4515 10854 4567 10906
rect 4579 10854 4631 10906
rect 7696 10854 7748 10906
rect 7760 10854 7812 10906
rect 7824 10854 7876 10906
rect 7888 10854 7940 10906
rect 7952 10854 8004 10906
rect 3700 10795 3752 10804
rect 3700 10761 3709 10795
rect 3709 10761 3743 10795
rect 3743 10761 3752 10795
rect 3700 10752 3752 10761
rect 9036 10795 9088 10804
rect 9036 10761 9045 10795
rect 9045 10761 9079 10795
rect 9079 10761 9088 10795
rect 9036 10752 9088 10761
rect 10140 10795 10192 10804
rect 10140 10761 10149 10795
rect 10149 10761 10183 10795
rect 10183 10761 10192 10795
rect 10140 10752 10192 10761
rect 7564 10727 7616 10736
rect 1768 10659 1820 10668
rect 1768 10625 1777 10659
rect 1777 10625 1811 10659
rect 1811 10625 1820 10659
rect 1768 10616 1820 10625
rect 7564 10693 7573 10727
rect 7573 10693 7607 10727
rect 7607 10693 7616 10727
rect 7564 10684 7616 10693
rect 3424 10616 3476 10668
rect 4068 10616 4120 10668
rect 6552 10659 6604 10668
rect 6552 10625 6561 10659
rect 6561 10625 6595 10659
rect 6595 10625 6604 10659
rect 6552 10616 6604 10625
rect 8668 10616 8720 10668
rect 1400 10591 1452 10600
rect 1400 10557 1409 10591
rect 1409 10557 1443 10591
rect 1443 10557 1452 10591
rect 1400 10548 1452 10557
rect 3056 10548 3108 10600
rect 5816 10548 5868 10600
rect 9772 10548 9824 10600
rect 9956 10548 10008 10600
rect 3148 10412 3200 10464
rect 5540 10412 5592 10464
rect 10324 10412 10376 10464
rect 2636 10310 2688 10362
rect 2700 10310 2752 10362
rect 2764 10310 2816 10362
rect 2828 10310 2880 10362
rect 2892 10310 2944 10362
rect 6010 10310 6062 10362
rect 6074 10310 6126 10362
rect 6138 10310 6190 10362
rect 6202 10310 6254 10362
rect 6266 10310 6318 10362
rect 9383 10310 9435 10362
rect 9447 10310 9499 10362
rect 9511 10310 9563 10362
rect 9575 10310 9627 10362
rect 9639 10310 9691 10362
rect 1492 10251 1544 10260
rect 1492 10217 1501 10251
rect 1501 10217 1535 10251
rect 1535 10217 1544 10251
rect 1492 10208 1544 10217
rect 3056 10208 3108 10260
rect 5632 10208 5684 10260
rect 8944 10251 8996 10260
rect 8944 10217 8953 10251
rect 8953 10217 8987 10251
rect 8987 10217 8996 10251
rect 8944 10208 8996 10217
rect 10048 10208 10100 10260
rect 4160 10140 4212 10192
rect 2872 10047 2924 10056
rect 2872 10013 2881 10047
rect 2881 10013 2915 10047
rect 2915 10013 2924 10047
rect 2872 10004 2924 10013
rect 3700 10072 3752 10124
rect 3148 10047 3200 10056
rect 3148 10013 3157 10047
rect 3157 10013 3191 10047
rect 3191 10013 3200 10047
rect 3148 10004 3200 10013
rect 4160 10047 4212 10056
rect 4160 10013 4169 10047
rect 4169 10013 4203 10047
rect 4203 10013 4212 10047
rect 4160 10004 4212 10013
rect 5540 10115 5592 10124
rect 5540 10081 5549 10115
rect 5549 10081 5583 10115
rect 5583 10081 5592 10115
rect 5540 10072 5592 10081
rect 7012 10072 7064 10124
rect 9772 10072 9824 10124
rect 3884 9936 3936 9988
rect 6828 10004 6880 10056
rect 9036 10004 9088 10056
rect 10324 10047 10376 10056
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 10324 10004 10376 10013
rect 5816 9868 5868 9920
rect 6552 9868 6604 9920
rect 6920 9868 6972 9920
rect 8392 9868 8444 9920
rect 4323 9766 4375 9818
rect 4387 9766 4439 9818
rect 4451 9766 4503 9818
rect 4515 9766 4567 9818
rect 4579 9766 4631 9818
rect 7696 9766 7748 9818
rect 7760 9766 7812 9818
rect 7824 9766 7876 9818
rect 7888 9766 7940 9818
rect 7952 9766 8004 9818
rect 3884 9707 3936 9716
rect 3884 9673 3893 9707
rect 3893 9673 3927 9707
rect 3927 9673 3936 9707
rect 3884 9664 3936 9673
rect 4160 9664 4212 9716
rect 6828 9664 6880 9716
rect 3424 9596 3476 9648
rect 7012 9596 7064 9648
rect 8208 9596 8260 9648
rect 8668 9596 8720 9648
rect 1400 9528 1452 9580
rect 4804 9571 4856 9580
rect 2412 9503 2464 9512
rect 2412 9469 2421 9503
rect 2421 9469 2455 9503
rect 2455 9469 2464 9503
rect 4804 9537 4813 9571
rect 4813 9537 4847 9571
rect 4847 9537 4856 9571
rect 4804 9528 4856 9537
rect 5356 9528 5408 9580
rect 2412 9460 2464 9469
rect 4896 9460 4948 9512
rect 6644 9460 6696 9512
rect 9220 9460 9272 9512
rect 9772 9460 9824 9512
rect 4252 9324 4304 9376
rect 9772 9324 9824 9376
rect 2636 9222 2688 9274
rect 2700 9222 2752 9274
rect 2764 9222 2816 9274
rect 2828 9222 2880 9274
rect 2892 9222 2944 9274
rect 6010 9222 6062 9274
rect 6074 9222 6126 9274
rect 6138 9222 6190 9274
rect 6202 9222 6254 9274
rect 6266 9222 6318 9274
rect 9383 9222 9435 9274
rect 9447 9222 9499 9274
rect 9511 9222 9563 9274
rect 9575 9222 9627 9274
rect 9639 9222 9691 9274
rect 4804 9120 4856 9172
rect 4160 8984 4212 9036
rect 8944 8984 8996 9036
rect 2044 8959 2096 8968
rect 2044 8925 2053 8959
rect 2053 8925 2087 8959
rect 2087 8925 2096 8959
rect 2044 8916 2096 8925
rect 4712 8959 4764 8968
rect 4712 8925 4721 8959
rect 4721 8925 4755 8959
rect 4755 8925 4764 8959
rect 4712 8916 4764 8925
rect 4804 8916 4856 8968
rect 5264 8916 5316 8968
rect 6644 8959 6696 8968
rect 6644 8925 6653 8959
rect 6653 8925 6687 8959
rect 6687 8925 6696 8959
rect 6644 8916 6696 8925
rect 8208 8916 8260 8968
rect 1676 8780 1728 8832
rect 5356 8780 5408 8832
rect 10232 8848 10284 8900
rect 8392 8823 8444 8832
rect 8392 8789 8401 8823
rect 8401 8789 8435 8823
rect 8435 8789 8444 8823
rect 8392 8780 8444 8789
rect 4323 8678 4375 8730
rect 4387 8678 4439 8730
rect 4451 8678 4503 8730
rect 4515 8678 4567 8730
rect 4579 8678 4631 8730
rect 7696 8678 7748 8730
rect 7760 8678 7812 8730
rect 7824 8678 7876 8730
rect 7888 8678 7940 8730
rect 7952 8678 8004 8730
rect 1400 8576 1452 8628
rect 3148 8576 3200 8628
rect 1676 8551 1728 8560
rect 1676 8517 1685 8551
rect 1685 8517 1719 8551
rect 1719 8517 1728 8551
rect 1676 8508 1728 8517
rect 3424 8508 3476 8560
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 2412 8372 2464 8424
rect 8760 8576 8812 8628
rect 9220 8619 9272 8628
rect 9220 8585 9229 8619
rect 9229 8585 9263 8619
rect 9263 8585 9272 8619
rect 9220 8576 9272 8585
rect 4252 8508 4304 8560
rect 3976 8372 4028 8424
rect 6552 8483 6604 8492
rect 6552 8449 6561 8483
rect 6561 8449 6595 8483
rect 6595 8449 6604 8483
rect 6552 8440 6604 8449
rect 7380 8508 7432 8560
rect 8024 8508 8076 8560
rect 8208 8508 8260 8560
rect 6920 8372 6972 8424
rect 5448 8304 5500 8356
rect 6644 8304 6696 8356
rect 2636 8134 2688 8186
rect 2700 8134 2752 8186
rect 2764 8134 2816 8186
rect 2828 8134 2880 8186
rect 2892 8134 2944 8186
rect 6010 8134 6062 8186
rect 6074 8134 6126 8186
rect 6138 8134 6190 8186
rect 6202 8134 6254 8186
rect 6266 8134 6318 8186
rect 9383 8134 9435 8186
rect 9447 8134 9499 8186
rect 9511 8134 9563 8186
rect 9575 8134 9627 8186
rect 9639 8134 9691 8186
rect 2044 8032 2096 8084
rect 4252 8032 4304 8084
rect 4712 8032 4764 8084
rect 8024 8075 8076 8084
rect 8024 8041 8033 8075
rect 8033 8041 8067 8075
rect 8067 8041 8076 8075
rect 8024 8032 8076 8041
rect 8944 8075 8996 8084
rect 8944 8041 8953 8075
rect 8953 8041 8987 8075
rect 8987 8041 8996 8075
rect 8944 8032 8996 8041
rect 8392 7964 8444 8016
rect 2044 7896 2096 7948
rect 2320 7896 2372 7948
rect 2412 7828 2464 7880
rect 5540 7871 5592 7880
rect 5540 7837 5549 7871
rect 5549 7837 5583 7871
rect 5583 7837 5592 7871
rect 6644 7896 6696 7948
rect 8760 7896 8812 7948
rect 5540 7828 5592 7837
rect 8024 7828 8076 7880
rect 3976 7760 4028 7812
rect 5264 7803 5316 7812
rect 5264 7769 5273 7803
rect 5273 7769 5307 7803
rect 5307 7769 5316 7803
rect 5264 7760 5316 7769
rect 6552 7803 6604 7812
rect 6552 7769 6561 7803
rect 6561 7769 6595 7803
rect 6595 7769 6604 7803
rect 6552 7760 6604 7769
rect 7012 7760 7064 7812
rect 5448 7692 5500 7744
rect 10416 7735 10468 7744
rect 10416 7701 10425 7735
rect 10425 7701 10459 7735
rect 10459 7701 10468 7735
rect 10416 7692 10468 7701
rect 4323 7590 4375 7642
rect 4387 7590 4439 7642
rect 4451 7590 4503 7642
rect 4515 7590 4567 7642
rect 4579 7590 4631 7642
rect 7696 7590 7748 7642
rect 7760 7590 7812 7642
rect 7824 7590 7876 7642
rect 7888 7590 7940 7642
rect 7952 7590 8004 7642
rect 3056 7488 3108 7540
rect 3976 7488 4028 7540
rect 4896 7531 4948 7540
rect 4896 7497 4905 7531
rect 4905 7497 4939 7531
rect 4939 7497 4948 7531
rect 4896 7488 4948 7497
rect 8024 7488 8076 7540
rect 4252 7420 4304 7472
rect 5080 7420 5132 7472
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 7564 7395 7616 7404
rect 7564 7361 7573 7395
rect 7573 7361 7607 7395
rect 7607 7361 7616 7395
rect 7564 7352 7616 7361
rect 4252 7327 4304 7336
rect 4252 7293 4261 7327
rect 4261 7293 4295 7327
rect 4295 7293 4304 7327
rect 4252 7284 4304 7293
rect 7380 7327 7432 7336
rect 7380 7293 7389 7327
rect 7389 7293 7423 7327
rect 7423 7293 7432 7327
rect 7380 7284 7432 7293
rect 8208 7420 8260 7472
rect 8944 7284 8996 7336
rect 10232 7327 10284 7336
rect 10232 7293 10241 7327
rect 10241 7293 10275 7327
rect 10275 7293 10284 7327
rect 10232 7284 10284 7293
rect 10508 7327 10560 7336
rect 10508 7293 10517 7327
rect 10517 7293 10551 7327
rect 10551 7293 10560 7327
rect 10508 7284 10560 7293
rect 5264 7216 5316 7268
rect 1400 7191 1452 7200
rect 1400 7157 1409 7191
rect 1409 7157 1443 7191
rect 1443 7157 1452 7191
rect 1400 7148 1452 7157
rect 2636 7046 2688 7098
rect 2700 7046 2752 7098
rect 2764 7046 2816 7098
rect 2828 7046 2880 7098
rect 2892 7046 2944 7098
rect 6010 7046 6062 7098
rect 6074 7046 6126 7098
rect 6138 7046 6190 7098
rect 6202 7046 6254 7098
rect 6266 7046 6318 7098
rect 9383 7046 9435 7098
rect 9447 7046 9499 7098
rect 9511 7046 9563 7098
rect 9575 7046 9627 7098
rect 9639 7046 9691 7098
rect 1492 6919 1544 6928
rect 1492 6885 1501 6919
rect 1501 6885 1535 6919
rect 1535 6885 1544 6919
rect 1492 6876 1544 6885
rect 7012 6876 7064 6928
rect 8208 6876 8260 6928
rect 6552 6808 6604 6860
rect 2412 6740 2464 6792
rect 3148 6740 3200 6792
rect 5540 6783 5592 6792
rect 5540 6749 5549 6783
rect 5549 6749 5583 6783
rect 5583 6749 5592 6783
rect 5540 6740 5592 6749
rect 8116 6740 8168 6792
rect 5816 6715 5868 6724
rect 5816 6681 5825 6715
rect 5825 6681 5859 6715
rect 5859 6681 5868 6715
rect 5816 6672 5868 6681
rect 9404 6740 9456 6792
rect 2964 6604 3016 6656
rect 3148 6604 3200 6656
rect 4068 6604 4120 6656
rect 10140 6672 10192 6724
rect 9864 6604 9916 6656
rect 4323 6502 4375 6554
rect 4387 6502 4439 6554
rect 4451 6502 4503 6554
rect 4515 6502 4567 6554
rect 4579 6502 4631 6554
rect 7696 6502 7748 6554
rect 7760 6502 7812 6554
rect 7824 6502 7876 6554
rect 7888 6502 7940 6554
rect 7952 6502 8004 6554
rect 5816 6443 5868 6452
rect 5816 6409 5825 6443
rect 5825 6409 5859 6443
rect 5859 6409 5868 6443
rect 5816 6400 5868 6409
rect 7564 6400 7616 6452
rect 10232 6400 10284 6452
rect 1400 6332 1452 6384
rect 3056 6332 3108 6384
rect 4068 6332 4120 6384
rect 8208 6332 8260 6384
rect 7104 6264 7156 6316
rect 2780 6196 2832 6248
rect 4344 6239 4396 6248
rect 4344 6205 4353 6239
rect 4353 6205 4387 6239
rect 4387 6205 4396 6239
rect 4344 6196 4396 6205
rect 8392 6239 8444 6248
rect 8392 6205 8401 6239
rect 8401 6205 8435 6239
rect 8435 6205 8444 6239
rect 8392 6196 8444 6205
rect 9036 6196 9088 6248
rect 9404 6196 9456 6248
rect 3424 6060 3476 6112
rect 2636 5958 2688 6010
rect 2700 5958 2752 6010
rect 2764 5958 2816 6010
rect 2828 5958 2880 6010
rect 2892 5958 2944 6010
rect 6010 5958 6062 6010
rect 6074 5958 6126 6010
rect 6138 5958 6190 6010
rect 6202 5958 6254 6010
rect 6266 5958 6318 6010
rect 9383 5958 9435 6010
rect 9447 5958 9499 6010
rect 9511 5958 9563 6010
rect 9575 5958 9627 6010
rect 9639 5958 9691 6010
rect 2504 5695 2556 5704
rect 2504 5661 2513 5695
rect 2513 5661 2547 5695
rect 2547 5661 2556 5695
rect 2504 5652 2556 5661
rect 3700 5652 3752 5704
rect 4160 5720 4212 5772
rect 4344 5720 4396 5772
rect 6920 5720 6972 5772
rect 8116 5763 8168 5772
rect 8116 5729 8125 5763
rect 8125 5729 8159 5763
rect 8159 5729 8168 5763
rect 8116 5720 8168 5729
rect 9036 5763 9088 5772
rect 9036 5729 9045 5763
rect 9045 5729 9079 5763
rect 9079 5729 9088 5763
rect 9036 5720 9088 5729
rect 3424 5584 3476 5636
rect 4804 5652 4856 5704
rect 7012 5652 7064 5704
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 8944 5652 8996 5704
rect 3148 5559 3200 5568
rect 3148 5525 3157 5559
rect 3157 5525 3191 5559
rect 3191 5525 3200 5559
rect 3148 5516 3200 5525
rect 7104 5516 7156 5568
rect 8116 5516 8168 5568
rect 9772 5516 9824 5568
rect 4323 5414 4375 5466
rect 4387 5414 4439 5466
rect 4451 5414 4503 5466
rect 4515 5414 4567 5466
rect 4579 5414 4631 5466
rect 7696 5414 7748 5466
rect 7760 5414 7812 5466
rect 7824 5414 7876 5466
rect 7888 5414 7940 5466
rect 7952 5414 8004 5466
rect 2320 5312 2372 5364
rect 3056 5312 3108 5364
rect 3424 5244 3476 5296
rect 4068 5312 4120 5364
rect 4160 5312 4212 5364
rect 5448 5244 5500 5296
rect 7012 5312 7064 5364
rect 8944 5312 8996 5364
rect 8116 5244 8168 5296
rect 8208 5244 8260 5296
rect 10140 5244 10192 5296
rect 10324 5244 10376 5296
rect 2872 5219 2924 5228
rect 2872 5185 2881 5219
rect 2881 5185 2915 5219
rect 2915 5185 2924 5219
rect 2872 5176 2924 5185
rect 5356 5219 5408 5228
rect 5356 5185 5365 5219
rect 5365 5185 5399 5219
rect 5399 5185 5408 5219
rect 5356 5176 5408 5185
rect 5632 5219 5684 5228
rect 5632 5185 5641 5219
rect 5641 5185 5675 5219
rect 5675 5185 5684 5219
rect 5632 5176 5684 5185
rect 5724 5176 5776 5228
rect 10508 5219 10560 5228
rect 10508 5185 10517 5219
rect 10517 5185 10551 5219
rect 10551 5185 10560 5219
rect 10508 5176 10560 5185
rect 6644 5108 6696 5160
rect 8392 5108 8444 5160
rect 4804 4972 4856 5024
rect 7196 4972 7248 5024
rect 2636 4870 2688 4922
rect 2700 4870 2752 4922
rect 2764 4870 2816 4922
rect 2828 4870 2880 4922
rect 2892 4870 2944 4922
rect 6010 4870 6062 4922
rect 6074 4870 6126 4922
rect 6138 4870 6190 4922
rect 6202 4870 6254 4922
rect 6266 4870 6318 4922
rect 9383 4870 9435 4922
rect 9447 4870 9499 4922
rect 9511 4870 9563 4922
rect 9575 4870 9627 4922
rect 9639 4870 9691 4922
rect 2504 4768 2556 4820
rect 3700 4768 3752 4820
rect 5632 4768 5684 4820
rect 3148 4700 3200 4752
rect 4896 4700 4948 4752
rect 4160 4632 4212 4684
rect 5172 4632 5224 4684
rect 2320 4496 2372 4548
rect 2964 4496 3016 4548
rect 5724 4564 5776 4616
rect 6368 4607 6420 4616
rect 6368 4573 6377 4607
rect 6377 4573 6411 4607
rect 6411 4573 6420 4607
rect 6368 4564 6420 4573
rect 5540 4496 5592 4548
rect 7472 4564 7524 4616
rect 8208 4632 8260 4684
rect 9312 4675 9364 4684
rect 9312 4641 9321 4675
rect 9321 4641 9355 4675
rect 9355 4641 9364 4675
rect 9312 4632 9364 4641
rect 10508 4607 10560 4616
rect 7196 4496 7248 4548
rect 10508 4573 10517 4607
rect 10517 4573 10551 4607
rect 10551 4573 10560 4607
rect 10508 4564 10560 4573
rect 8208 4496 8260 4548
rect 4252 4471 4304 4480
rect 4252 4437 4261 4471
rect 4261 4437 4295 4471
rect 4295 4437 4304 4471
rect 4252 4428 4304 4437
rect 4988 4471 5040 4480
rect 4988 4437 4997 4471
rect 4997 4437 5031 4471
rect 5031 4437 5040 4471
rect 4988 4428 5040 4437
rect 5264 4428 5316 4480
rect 6920 4428 6972 4480
rect 4323 4326 4375 4378
rect 4387 4326 4439 4378
rect 4451 4326 4503 4378
rect 4515 4326 4567 4378
rect 4579 4326 4631 4378
rect 7696 4326 7748 4378
rect 7760 4326 7812 4378
rect 7824 4326 7876 4378
rect 7888 4326 7940 4378
rect 7952 4326 8004 4378
rect 5356 4224 5408 4276
rect 5540 4224 5592 4276
rect 7472 4224 7524 4276
rect 10324 4224 10376 4276
rect 4160 4156 4212 4208
rect 9312 4156 9364 4208
rect 2136 4131 2188 4140
rect 2136 4097 2145 4131
rect 2145 4097 2179 4131
rect 2179 4097 2188 4131
rect 2136 4088 2188 4097
rect 4988 4088 5040 4140
rect 5448 4088 5500 4140
rect 2228 4020 2280 4072
rect 4344 4020 4396 4072
rect 5080 4020 5132 4072
rect 6368 4020 6420 4072
rect 7196 4020 7248 4072
rect 2044 3952 2096 4004
rect 5172 3952 5224 4004
rect 1492 3927 1544 3936
rect 1492 3893 1501 3927
rect 1501 3893 1535 3927
rect 1535 3893 1544 3927
rect 1492 3884 1544 3893
rect 2504 3884 2556 3936
rect 3884 3884 3936 3936
rect 6368 3927 6420 3936
rect 6368 3893 6377 3927
rect 6377 3893 6411 3927
rect 6411 3893 6420 3927
rect 6368 3884 6420 3893
rect 6644 3884 6696 3936
rect 9036 4063 9088 4072
rect 9036 4029 9045 4063
rect 9045 4029 9079 4063
rect 9079 4029 9088 4063
rect 9036 4020 9088 4029
rect 2636 3782 2688 3834
rect 2700 3782 2752 3834
rect 2764 3782 2816 3834
rect 2828 3782 2880 3834
rect 2892 3782 2944 3834
rect 6010 3782 6062 3834
rect 6074 3782 6126 3834
rect 6138 3782 6190 3834
rect 6202 3782 6254 3834
rect 6266 3782 6318 3834
rect 9383 3782 9435 3834
rect 9447 3782 9499 3834
rect 9511 3782 9563 3834
rect 9575 3782 9627 3834
rect 9639 3782 9691 3834
rect 2136 3680 2188 3732
rect 5724 3680 5776 3732
rect 2044 3587 2096 3596
rect 2044 3553 2053 3587
rect 2053 3553 2087 3587
rect 2087 3553 2096 3587
rect 2044 3544 2096 3553
rect 2412 3544 2464 3596
rect 2964 3544 3016 3596
rect 4068 3587 4120 3596
rect 4068 3553 4077 3587
rect 4077 3553 4111 3587
rect 4111 3553 4120 3587
rect 4068 3544 4120 3553
rect 4804 3544 4856 3596
rect 6644 3519 6696 3528
rect 6644 3485 6653 3519
rect 6653 3485 6687 3519
rect 6687 3485 6696 3519
rect 6644 3476 6696 3485
rect 8024 3476 8076 3528
rect 9772 3612 9824 3664
rect 9864 3544 9916 3596
rect 2228 3383 2280 3392
rect 2228 3349 2237 3383
rect 2237 3349 2271 3383
rect 2271 3349 2280 3383
rect 2228 3340 2280 3349
rect 4160 3340 4212 3392
rect 9956 3476 10008 3528
rect 4323 3238 4375 3290
rect 4387 3238 4439 3290
rect 4451 3238 4503 3290
rect 4515 3238 4567 3290
rect 4579 3238 4631 3290
rect 7696 3238 7748 3290
rect 7760 3238 7812 3290
rect 7824 3238 7876 3290
rect 7888 3238 7940 3290
rect 7952 3238 8004 3290
rect 2228 3136 2280 3188
rect 2504 3136 2556 3188
rect 5264 3136 5316 3188
rect 2320 3068 2372 3120
rect 2964 3068 3016 3120
rect 3884 3111 3936 3120
rect 3884 3077 3893 3111
rect 3893 3077 3927 3111
rect 3927 3077 3936 3111
rect 3884 3068 3936 3077
rect 4160 3068 4212 3120
rect 9036 3136 9088 3188
rect 6368 3068 6420 3120
rect 8024 3068 8076 3120
rect 6644 3000 6696 3052
rect 6460 2796 6512 2848
rect 2636 2694 2688 2746
rect 2700 2694 2752 2746
rect 2764 2694 2816 2746
rect 2828 2694 2880 2746
rect 2892 2694 2944 2746
rect 6010 2694 6062 2746
rect 6074 2694 6126 2746
rect 6138 2694 6190 2746
rect 6202 2694 6254 2746
rect 6266 2694 6318 2746
rect 9383 2694 9435 2746
rect 9447 2694 9499 2746
rect 9511 2694 9563 2746
rect 9575 2694 9627 2746
rect 9639 2694 9691 2746
rect 8208 2592 8260 2644
rect 4252 2524 4304 2576
rect 4160 2499 4212 2508
rect 4160 2465 4169 2499
rect 4169 2465 4203 2499
rect 4203 2465 4212 2499
rect 6644 2499 6696 2508
rect 4160 2456 4212 2465
rect 6644 2465 6653 2499
rect 6653 2465 6687 2499
rect 6687 2465 6696 2499
rect 6644 2456 6696 2465
rect 6920 2499 6972 2508
rect 6920 2465 6929 2499
rect 6929 2465 6963 2499
rect 6963 2465 6972 2499
rect 6920 2456 6972 2465
rect 3240 2388 3292 2440
rect 8024 2388 8076 2440
rect 9956 2388 10008 2440
rect 20 2320 72 2372
rect 9680 2295 9732 2304
rect 9680 2261 9689 2295
rect 9689 2261 9723 2295
rect 9723 2261 9732 2295
rect 9680 2252 9732 2261
rect 10416 2295 10468 2304
rect 10416 2261 10425 2295
rect 10425 2261 10459 2295
rect 10459 2261 10468 2295
rect 10416 2252 10468 2261
rect 4323 2150 4375 2202
rect 4387 2150 4439 2202
rect 4451 2150 4503 2202
rect 4515 2150 4567 2202
rect 4579 2150 4631 2202
rect 7696 2150 7748 2202
rect 7760 2150 7812 2202
rect 7824 2150 7876 2202
rect 7888 2150 7940 2202
rect 7952 2150 8004 2202
<< metal2 >>
rect 2594 13818 2650 14473
rect 2594 13790 2728 13818
rect 1490 13696 1546 13705
rect 2594 13673 2650 13790
rect 1490 13631 1546 13640
rect 1504 11898 1532 13631
rect 1492 11892 1544 11898
rect 1492 11834 1544 11840
rect 2700 11762 2728 13790
rect 5814 13673 5870 14473
rect 9034 13818 9090 14473
rect 9034 13790 9260 13818
rect 9034 13673 9090 13790
rect 4323 11996 4631 12016
rect 4323 11994 4329 11996
rect 4385 11994 4409 11996
rect 4465 11994 4489 11996
rect 4545 11994 4569 11996
rect 4625 11994 4631 11996
rect 4385 11942 4387 11994
rect 4567 11942 4569 11994
rect 4323 11940 4329 11942
rect 4385 11940 4409 11942
rect 4465 11940 4489 11942
rect 4545 11940 4569 11942
rect 4625 11940 4631 11942
rect 4323 11920 4631 11940
rect 5828 11898 5856 13673
rect 7696 11996 8004 12016
rect 7696 11994 7702 11996
rect 7758 11994 7782 11996
rect 7838 11994 7862 11996
rect 7918 11994 7942 11996
rect 7998 11994 8004 11996
rect 7758 11942 7760 11994
rect 7940 11942 7942 11994
rect 7696 11940 7702 11942
rect 7758 11940 7782 11942
rect 7838 11940 7862 11942
rect 7918 11940 7942 11942
rect 7998 11940 8004 11942
rect 7696 11920 8004 11940
rect 9232 11898 9260 13790
rect 12254 13673 12310 14473
rect 12268 11898 12296 13673
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2688 11756 2740 11762
rect 2688 11698 2740 11704
rect 5724 11756 5776 11762
rect 5724 11698 5776 11704
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1780 10674 1808 11086
rect 1768 10668 1820 10674
rect 1768 10610 1820 10616
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1412 9586 1440 10542
rect 1490 10296 1546 10305
rect 1490 10231 1492 10240
rect 1544 10231 1546 10240
rect 1492 10202 1544 10208
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1412 8634 1440 9522
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1400 8628 1452 8634
rect 1400 8570 1452 8576
rect 1412 8498 1440 8570
rect 1688 8566 1716 8774
rect 1676 8560 1728 8566
rect 1676 8502 1728 8508
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 2056 8090 2084 8910
rect 2424 8514 2452 9454
rect 2332 8486 2452 8514
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 2332 7954 2360 8486
rect 2412 8424 2464 8430
rect 2412 8366 2464 8372
rect 2044 7948 2096 7954
rect 2044 7890 2096 7896
rect 2320 7948 2372 7954
rect 2320 7890 2372 7896
rect 1400 7200 1452 7206
rect 1400 7142 1452 7148
rect 1412 6390 1440 7142
rect 1492 6928 1544 6934
rect 1490 6896 1492 6905
rect 1544 6896 1546 6905
rect 1490 6831 1546 6840
rect 1400 6384 1452 6390
rect 1400 6326 1452 6332
rect 2056 4010 2084 7890
rect 2424 7886 2452 8366
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2424 6798 2452 7822
rect 2412 6792 2464 6798
rect 2412 6734 2464 6740
rect 2516 5710 2544 11698
rect 3700 11620 3752 11626
rect 3700 11562 3752 11568
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2636 11452 2944 11472
rect 2636 11450 2642 11452
rect 2698 11450 2722 11452
rect 2778 11450 2802 11452
rect 2858 11450 2882 11452
rect 2938 11450 2944 11452
rect 2698 11398 2700 11450
rect 2880 11398 2882 11450
rect 2636 11396 2642 11398
rect 2698 11396 2722 11398
rect 2778 11396 2802 11398
rect 2858 11396 2882 11398
rect 2938 11396 2944 11398
rect 2636 11376 2944 11396
rect 2636 10364 2944 10384
rect 2636 10362 2642 10364
rect 2698 10362 2722 10364
rect 2778 10362 2802 10364
rect 2858 10362 2882 10364
rect 2938 10362 2944 10364
rect 2698 10310 2700 10362
rect 2880 10310 2882 10362
rect 2636 10308 2642 10310
rect 2698 10308 2722 10310
rect 2778 10308 2802 10310
rect 2858 10308 2882 10310
rect 2938 10308 2944 10310
rect 2636 10288 2944 10308
rect 2976 10146 3004 11494
rect 3712 10810 3740 11562
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 3700 10804 3752 10810
rect 3700 10746 3752 10752
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 3068 10266 3096 10542
rect 3148 10464 3200 10470
rect 3148 10406 3200 10412
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 2884 10118 3004 10146
rect 2884 10062 2912 10118
rect 3160 10062 3188 10406
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3436 9654 3464 10610
rect 3712 10130 3740 10746
rect 4080 10674 4108 11018
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 4172 10198 4200 10950
rect 4323 10908 4631 10928
rect 4323 10906 4329 10908
rect 4385 10906 4409 10908
rect 4465 10906 4489 10908
rect 4545 10906 4569 10908
rect 4625 10906 4631 10908
rect 4385 10854 4387 10906
rect 4567 10854 4569 10906
rect 4323 10852 4329 10854
rect 4385 10852 4409 10854
rect 4465 10852 4489 10854
rect 4545 10852 4569 10854
rect 4625 10852 4631 10854
rect 4323 10832 4631 10852
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 4160 10192 4212 10198
rect 4160 10134 4212 10140
rect 5552 10130 5580 10406
rect 5644 10266 5672 11018
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 3884 9988 3936 9994
rect 3884 9930 3936 9936
rect 3896 9722 3924 9930
rect 4172 9722 4200 9998
rect 4323 9820 4631 9840
rect 4323 9818 4329 9820
rect 4385 9818 4409 9820
rect 4465 9818 4489 9820
rect 4545 9818 4569 9820
rect 4625 9818 4631 9820
rect 4385 9766 4387 9818
rect 4567 9766 4569 9818
rect 4323 9764 4329 9766
rect 4385 9764 4409 9766
rect 4465 9764 4489 9766
rect 4545 9764 4569 9766
rect 4625 9764 4631 9766
rect 4323 9744 4631 9764
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 4160 9716 4212 9722
rect 4160 9658 4212 9664
rect 3424 9648 3476 9654
rect 3424 9590 3476 9596
rect 2636 9276 2944 9296
rect 2636 9274 2642 9276
rect 2698 9274 2722 9276
rect 2778 9274 2802 9276
rect 2858 9274 2882 9276
rect 2938 9274 2944 9276
rect 2698 9222 2700 9274
rect 2880 9222 2882 9274
rect 2636 9220 2642 9222
rect 2698 9220 2722 9222
rect 2778 9220 2802 9222
rect 2858 9220 2882 9222
rect 2938 9220 2944 9222
rect 2636 9200 2944 9220
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 2636 8188 2944 8208
rect 2636 8186 2642 8188
rect 2698 8186 2722 8188
rect 2778 8186 2802 8188
rect 2858 8186 2882 8188
rect 2938 8186 2944 8188
rect 2698 8134 2700 8186
rect 2880 8134 2882 8186
rect 2636 8132 2642 8134
rect 2698 8132 2722 8134
rect 2778 8132 2802 8134
rect 2858 8132 2882 8134
rect 2938 8132 2944 8134
rect 2636 8112 2944 8132
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 2636 7100 2944 7120
rect 2636 7098 2642 7100
rect 2698 7098 2722 7100
rect 2778 7098 2802 7100
rect 2858 7098 2882 7100
rect 2938 7098 2944 7100
rect 2698 7046 2700 7098
rect 2880 7046 2882 7098
rect 2636 7044 2642 7046
rect 2698 7044 2722 7046
rect 2778 7044 2802 7046
rect 2858 7044 2882 7046
rect 2938 7044 2944 7046
rect 2636 7024 2944 7044
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2780 6248 2832 6254
rect 2976 6202 3004 6598
rect 3068 6390 3096 7482
rect 3160 7410 3188 8570
rect 3436 8566 3464 9590
rect 4172 9042 4200 9658
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 4264 8566 4292 9318
rect 4816 9178 4844 9522
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4323 8732 4631 8752
rect 4323 8730 4329 8732
rect 4385 8730 4409 8732
rect 4465 8730 4489 8732
rect 4545 8730 4569 8732
rect 4625 8730 4631 8732
rect 4385 8678 4387 8730
rect 4567 8678 4569 8730
rect 4323 8676 4329 8678
rect 4385 8676 4409 8678
rect 4465 8676 4489 8678
rect 4545 8676 4569 8678
rect 4625 8676 4631 8678
rect 4323 8656 4631 8676
rect 3424 8560 3476 8566
rect 3424 8502 3476 8508
rect 4252 8560 4304 8566
rect 4252 8502 4304 8508
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 3988 7818 4016 8366
rect 4724 8090 4752 8910
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 3988 7546 4016 7754
rect 3976 7540 4028 7546
rect 3976 7482 4028 7488
rect 4264 7478 4292 8026
rect 4323 7644 4631 7664
rect 4323 7642 4329 7644
rect 4385 7642 4409 7644
rect 4465 7642 4489 7644
rect 4545 7642 4569 7644
rect 4625 7642 4631 7644
rect 4385 7590 4387 7642
rect 4567 7590 4569 7642
rect 4323 7588 4329 7590
rect 4385 7588 4409 7590
rect 4465 7588 4489 7590
rect 4545 7588 4569 7590
rect 4625 7588 4631 7590
rect 4323 7568 4631 7588
rect 4252 7472 4304 7478
rect 4252 7414 4304 7420
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3160 6798 3188 7346
rect 4264 7342 4292 7414
rect 4252 7336 4304 7342
rect 4252 7278 4304 7284
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3160 6662 3188 6734
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 4080 6390 4108 6598
rect 4323 6556 4631 6576
rect 4323 6554 4329 6556
rect 4385 6554 4409 6556
rect 4465 6554 4489 6556
rect 4545 6554 4569 6556
rect 4625 6554 4631 6556
rect 4385 6502 4387 6554
rect 4567 6502 4569 6554
rect 4323 6500 4329 6502
rect 4385 6500 4409 6502
rect 4465 6500 4489 6502
rect 4545 6500 4569 6502
rect 4625 6500 4631 6502
rect 4323 6480 4631 6500
rect 3056 6384 3108 6390
rect 3056 6326 3108 6332
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 2832 6196 3004 6202
rect 2780 6190 3004 6196
rect 2792 6174 3004 6190
rect 2636 6012 2944 6032
rect 2636 6010 2642 6012
rect 2698 6010 2722 6012
rect 2778 6010 2802 6012
rect 2858 6010 2882 6012
rect 2938 6010 2944 6012
rect 2698 5958 2700 6010
rect 2880 5958 2882 6010
rect 2636 5956 2642 5958
rect 2698 5956 2722 5958
rect 2778 5956 2802 5958
rect 2858 5956 2882 5958
rect 2938 5956 2944 5958
rect 2636 5936 2944 5956
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2320 5364 2372 5370
rect 2320 5306 2372 5312
rect 2332 4554 2360 5306
rect 2516 4826 2544 5646
rect 2976 5250 3004 6174
rect 3068 5370 3096 6326
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3436 5642 3464 6054
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3424 5636 3476 5642
rect 3424 5578 3476 5584
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 2884 5234 3004 5250
rect 2872 5228 3004 5234
rect 2924 5222 3004 5228
rect 2872 5170 2924 5176
rect 2636 4924 2944 4944
rect 2636 4922 2642 4924
rect 2698 4922 2722 4924
rect 2778 4922 2802 4924
rect 2858 4922 2882 4924
rect 2938 4922 2944 4924
rect 2698 4870 2700 4922
rect 2880 4870 2882 4922
rect 2636 4868 2642 4870
rect 2698 4868 2722 4870
rect 2778 4868 2802 4870
rect 2858 4868 2882 4870
rect 2938 4868 2944 4870
rect 2636 4848 2944 4868
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2320 4548 2372 4554
rect 2320 4490 2372 4496
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2044 4004 2096 4010
rect 2044 3946 2096 3952
rect 1492 3936 1544 3942
rect 1492 3878 1544 3884
rect 1504 3505 1532 3878
rect 2056 3602 2084 3946
rect 2148 3738 2176 4082
rect 2228 4072 2280 4078
rect 2228 4014 2280 4020
rect 2136 3732 2188 3738
rect 2136 3674 2188 3680
rect 2044 3596 2096 3602
rect 2044 3538 2096 3544
rect 1490 3496 1546 3505
rect 1490 3431 1546 3440
rect 2240 3398 2268 4014
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 2240 3194 2268 3334
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2332 3126 2360 4490
rect 2516 4026 2544 4762
rect 2976 4554 3004 5222
rect 3160 4758 3188 5510
rect 3436 5302 3464 5578
rect 3424 5296 3476 5302
rect 3424 5238 3476 5244
rect 3712 4826 3740 5646
rect 4080 5370 4108 6326
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 4356 5778 4384 6190
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4172 5370 4200 5714
rect 4816 5710 4844 8910
rect 4908 7546 4936 9454
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5276 7818 5304 8910
rect 5368 8838 5396 9522
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5368 8378 5396 8774
rect 5368 8362 5488 8378
rect 5368 8356 5500 8362
rect 5368 8350 5448 8356
rect 5448 8298 5500 8304
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 5080 7472 5132 7478
rect 5080 7414 5132 7420
rect 4804 5704 4856 5710
rect 4856 5664 4936 5692
rect 4804 5646 4856 5652
rect 4323 5468 4631 5488
rect 4323 5466 4329 5468
rect 4385 5466 4409 5468
rect 4465 5466 4489 5468
rect 4545 5466 4569 5468
rect 4625 5466 4631 5468
rect 4385 5414 4387 5466
rect 4567 5414 4569 5466
rect 4323 5412 4329 5414
rect 4385 5412 4409 5414
rect 4465 5412 4489 5414
rect 4545 5412 4569 5414
rect 4625 5412 4631 5414
rect 4323 5392 4631 5412
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3148 4752 3200 4758
rect 3148 4694 3200 4700
rect 2964 4548 3016 4554
rect 2964 4490 3016 4496
rect 2424 3998 2544 4026
rect 2424 3602 2452 3998
rect 2504 3936 2556 3942
rect 2504 3878 2556 3884
rect 2412 3596 2464 3602
rect 2412 3538 2464 3544
rect 2516 3194 2544 3878
rect 2636 3836 2944 3856
rect 2636 3834 2642 3836
rect 2698 3834 2722 3836
rect 2778 3834 2802 3836
rect 2858 3834 2882 3836
rect 2938 3834 2944 3836
rect 2698 3782 2700 3834
rect 2880 3782 2882 3834
rect 2636 3780 2642 3782
rect 2698 3780 2722 3782
rect 2778 3780 2802 3782
rect 2858 3780 2882 3782
rect 2938 3780 2944 3782
rect 2636 3760 2944 3780
rect 2976 3602 3004 4490
rect 4080 4162 4108 5306
rect 4172 4690 4200 5306
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4172 4214 4200 4245
rect 4160 4208 4212 4214
rect 4080 4156 4160 4162
rect 4080 4150 4212 4156
rect 4080 4134 4200 4150
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 2964 3596 3016 3602
rect 2964 3538 3016 3544
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2976 3126 3004 3538
rect 3896 3126 3924 3878
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 2320 3120 2372 3126
rect 2320 3062 2372 3068
rect 2964 3120 3016 3126
rect 2964 3062 3016 3068
rect 3884 3120 3936 3126
rect 3884 3062 3936 3068
rect 4080 2802 4108 3538
rect 4172 3398 4200 4134
rect 4264 4060 4292 4422
rect 4323 4380 4631 4400
rect 4323 4378 4329 4380
rect 4385 4378 4409 4380
rect 4465 4378 4489 4380
rect 4545 4378 4569 4380
rect 4625 4378 4631 4380
rect 4385 4326 4387 4378
rect 4567 4326 4569 4378
rect 4323 4324 4329 4326
rect 4385 4324 4409 4326
rect 4465 4324 4489 4326
rect 4545 4324 4569 4326
rect 4625 4324 4631 4326
rect 4323 4304 4631 4324
rect 4344 4072 4396 4078
rect 4264 4032 4344 4060
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 4172 3126 4200 3334
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 4080 2774 4200 2802
rect 2636 2748 2944 2768
rect 2636 2746 2642 2748
rect 2698 2746 2722 2748
rect 2778 2746 2802 2748
rect 2858 2746 2882 2748
rect 2938 2746 2944 2748
rect 2698 2694 2700 2746
rect 2880 2694 2882 2746
rect 2636 2692 2642 2694
rect 2698 2692 2722 2694
rect 2778 2692 2802 2694
rect 2858 2692 2882 2694
rect 2938 2692 2944 2694
rect 2636 2672 2944 2692
rect 4172 2514 4200 2774
rect 4264 2582 4292 4032
rect 4344 4014 4396 4020
rect 4816 3602 4844 4966
rect 4908 4758 4936 5664
rect 4896 4752 4948 4758
rect 4896 4694 4948 4700
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 5000 4146 5028 4422
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 5092 4078 5120 7414
rect 5276 7274 5304 7754
rect 5460 7750 5488 8298
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5264 7268 5316 7274
rect 5264 7210 5316 7216
rect 5552 6798 5580 7822
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5448 5296 5500 5302
rect 5448 5238 5500 5244
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 5184 4010 5212 4626
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 4323 3292 4631 3312
rect 4323 3290 4329 3292
rect 4385 3290 4409 3292
rect 4465 3290 4489 3292
rect 4545 3290 4569 3292
rect 4625 3290 4631 3292
rect 4385 3238 4387 3290
rect 4567 3238 4569 3290
rect 4323 3236 4329 3238
rect 4385 3236 4409 3238
rect 4465 3236 4489 3238
rect 4545 3236 4569 3238
rect 4625 3236 4631 3238
rect 4323 3216 4631 3236
rect 5276 3194 5304 4422
rect 5368 4282 5396 5170
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5460 4146 5488 5238
rect 5736 5234 5764 11698
rect 6552 11552 6604 11558
rect 6552 11494 6604 11500
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 6010 11452 6318 11472
rect 6010 11450 6016 11452
rect 6072 11450 6096 11452
rect 6152 11450 6176 11452
rect 6232 11450 6256 11452
rect 6312 11450 6318 11452
rect 6072 11398 6074 11450
rect 6254 11398 6256 11450
rect 6010 11396 6016 11398
rect 6072 11396 6096 11398
rect 6152 11396 6176 11398
rect 6232 11396 6256 11398
rect 6312 11396 6318 11398
rect 6010 11376 6318 11396
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 5920 10690 5948 11086
rect 5828 10662 5948 10690
rect 6564 10674 6592 11494
rect 7576 10742 7604 11494
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 7696 10908 8004 10928
rect 7696 10906 7702 10908
rect 7758 10906 7782 10908
rect 7838 10906 7862 10908
rect 7918 10906 7942 10908
rect 7998 10906 8004 10908
rect 7758 10854 7760 10906
rect 7940 10854 7942 10906
rect 7696 10852 7702 10854
rect 7758 10852 7782 10854
rect 7838 10852 7862 10854
rect 7918 10852 7942 10854
rect 7998 10852 8004 10854
rect 7696 10832 8004 10852
rect 7564 10736 7616 10742
rect 7564 10678 7616 10684
rect 8680 10674 8708 11018
rect 6552 10668 6604 10674
rect 5828 10606 5856 10662
rect 6552 10610 6604 10616
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5828 9926 5856 10542
rect 6010 10364 6318 10384
rect 6010 10362 6016 10364
rect 6072 10362 6096 10364
rect 6152 10362 6176 10364
rect 6232 10362 6256 10364
rect 6312 10362 6318 10364
rect 6072 10310 6074 10362
rect 6254 10310 6256 10362
rect 6010 10308 6016 10310
rect 6072 10308 6096 10310
rect 6152 10308 6176 10310
rect 6232 10308 6256 10310
rect 6312 10308 6318 10310
rect 6010 10288 6318 10308
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 5816 9920 5868 9926
rect 5816 9862 5868 9868
rect 6552 9920 6604 9926
rect 6604 9880 6684 9908
rect 6552 9862 6604 9868
rect 6656 9518 6684 9880
rect 6840 9722 6868 9998
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6010 9276 6318 9296
rect 6010 9274 6016 9276
rect 6072 9274 6096 9276
rect 6152 9274 6176 9276
rect 6232 9274 6256 9276
rect 6312 9274 6318 9276
rect 6072 9222 6074 9274
rect 6254 9222 6256 9274
rect 6010 9220 6016 9222
rect 6072 9220 6096 9222
rect 6152 9220 6176 9222
rect 6232 9220 6256 9222
rect 6312 9220 6318 9222
rect 6010 9200 6318 9220
rect 6656 8974 6684 9454
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6010 8188 6318 8208
rect 6010 8186 6016 8188
rect 6072 8186 6096 8188
rect 6152 8186 6176 8188
rect 6232 8186 6256 8188
rect 6312 8186 6318 8188
rect 6072 8134 6074 8186
rect 6254 8134 6256 8186
rect 6010 8132 6016 8134
rect 6072 8132 6096 8134
rect 6152 8132 6176 8134
rect 6232 8132 6256 8134
rect 6312 8132 6318 8134
rect 6010 8112 6318 8132
rect 6564 7818 6592 8434
rect 6656 8362 6684 8910
rect 6932 8430 6960 9862
rect 7024 9654 7052 10066
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 7696 9820 8004 9840
rect 7696 9818 7702 9820
rect 7758 9818 7782 9820
rect 7838 9818 7862 9820
rect 7918 9818 7942 9820
rect 7998 9818 8004 9820
rect 7758 9766 7760 9818
rect 7940 9766 7942 9818
rect 7696 9764 7702 9766
rect 7758 9764 7782 9766
rect 7838 9764 7862 9766
rect 7918 9764 7942 9766
rect 7998 9764 8004 9766
rect 7696 9744 8004 9764
rect 7012 9648 7064 9654
rect 7012 9590 7064 9596
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 8220 8974 8248 9590
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 7696 8732 8004 8752
rect 7696 8730 7702 8732
rect 7758 8730 7782 8732
rect 7838 8730 7862 8732
rect 7918 8730 7942 8732
rect 7998 8730 8004 8732
rect 7758 8678 7760 8730
rect 7940 8678 7942 8730
rect 7696 8676 7702 8678
rect 7758 8676 7782 8678
rect 7838 8676 7862 8678
rect 7918 8676 7942 8678
rect 7998 8676 8004 8678
rect 7696 8656 8004 8676
rect 8220 8566 8248 8910
rect 8404 8838 8432 9862
rect 8680 9654 8708 10610
rect 8956 10266 8984 11698
rect 9048 10810 9076 11698
rect 9383 11452 9691 11472
rect 9383 11450 9389 11452
rect 9445 11450 9469 11452
rect 9525 11450 9549 11452
rect 9605 11450 9629 11452
rect 9685 11450 9691 11452
rect 9445 11398 9447 11450
rect 9627 11398 9629 11450
rect 9383 11396 9389 11398
rect 9445 11396 9469 11398
rect 9525 11396 9549 11398
rect 9605 11396 9629 11398
rect 9685 11396 9691 11398
rect 9383 11376 9691 11396
rect 10152 11218 10180 11698
rect 10416 11280 10468 11286
rect 10416 11222 10468 11228
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 9036 10804 9088 10810
rect 9036 10746 9088 10752
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 9048 10062 9076 10746
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9383 10364 9691 10384
rect 9383 10362 9389 10364
rect 9445 10362 9469 10364
rect 9525 10362 9549 10364
rect 9605 10362 9629 10364
rect 9685 10362 9691 10364
rect 9445 10310 9447 10362
rect 9627 10310 9629 10362
rect 9383 10308 9389 10310
rect 9445 10308 9469 10310
rect 9525 10308 9549 10310
rect 9605 10308 9629 10310
rect 9685 10308 9691 10310
rect 9383 10288 9691 10308
rect 9784 10130 9812 10542
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 8668 9648 8720 9654
rect 8668 9590 8720 9596
rect 9784 9518 9812 10066
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 7380 8560 7432 8566
rect 7380 8502 7432 8508
rect 8024 8560 8076 8566
rect 8024 8502 8076 8508
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6656 7954 6684 8298
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6552 7812 6604 7818
rect 6552 7754 6604 7760
rect 6010 7100 6318 7120
rect 6010 7098 6016 7100
rect 6072 7098 6096 7100
rect 6152 7098 6176 7100
rect 6232 7098 6256 7100
rect 6312 7098 6318 7100
rect 6072 7046 6074 7098
rect 6254 7046 6256 7098
rect 6010 7044 6016 7046
rect 6072 7044 6096 7046
rect 6152 7044 6176 7046
rect 6232 7044 6256 7046
rect 6312 7044 6318 7046
rect 6010 7024 6318 7044
rect 6564 6866 6592 7754
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 5828 6458 5856 6666
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 6010 6012 6318 6032
rect 6010 6010 6016 6012
rect 6072 6010 6096 6012
rect 6152 6010 6176 6012
rect 6232 6010 6256 6012
rect 6312 6010 6318 6012
rect 6072 5958 6074 6010
rect 6254 5958 6256 6010
rect 6010 5956 6016 5958
rect 6072 5956 6096 5958
rect 6152 5956 6176 5958
rect 6232 5956 6256 5958
rect 6312 5956 6318 5958
rect 6010 5936 6318 5956
rect 6932 5778 6960 8366
rect 7012 7812 7064 7818
rect 7012 7754 7064 7760
rect 7024 6934 7052 7754
rect 7392 7342 7420 8502
rect 8036 8090 8064 8502
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 7696 7644 8004 7664
rect 7696 7642 7702 7644
rect 7758 7642 7782 7644
rect 7838 7642 7862 7644
rect 7918 7642 7942 7644
rect 7998 7642 8004 7644
rect 7758 7590 7760 7642
rect 7940 7590 7942 7642
rect 7696 7588 7702 7590
rect 7758 7588 7782 7590
rect 7838 7588 7862 7590
rect 7918 7588 7942 7590
rect 7998 7588 8004 7590
rect 7696 7568 8004 7588
rect 8036 7546 8064 7822
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 8220 7478 8248 8502
rect 8404 8022 8432 8774
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8392 8016 8444 8022
rect 8392 7958 8444 7964
rect 8772 7954 8800 8570
rect 8956 8090 8984 8978
rect 9232 8634 9260 9454
rect 9784 9382 9812 9454
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9383 9276 9691 9296
rect 9383 9274 9389 9276
rect 9445 9274 9469 9276
rect 9525 9274 9549 9276
rect 9605 9274 9629 9276
rect 9685 9274 9691 9276
rect 9445 9222 9447 9274
rect 9627 9222 9629 9274
rect 9383 9220 9389 9222
rect 9445 9220 9469 9222
rect 9525 9220 9549 9222
rect 9605 9220 9629 9222
rect 9685 9220 9691 9222
rect 9383 9200 9691 9220
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9383 8188 9691 8208
rect 9383 8186 9389 8188
rect 9445 8186 9469 8188
rect 9525 8186 9549 8188
rect 9605 8186 9629 8188
rect 9685 8186 9691 8188
rect 9445 8134 9447 8186
rect 9627 8134 9629 8186
rect 9383 8132 9389 8134
rect 9445 8132 9469 8134
rect 9525 8132 9549 8134
rect 9605 8132 9629 8134
rect 9685 8132 9691 8134
rect 9383 8112 9691 8132
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8208 7472 8260 7478
rect 8208 7414 8260 7420
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7012 6928 7064 6934
rect 7012 6870 7064 6876
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 7024 5710 7052 6870
rect 7576 6458 7604 7346
rect 8220 6934 8248 7414
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 7696 6556 8004 6576
rect 7696 6554 7702 6556
rect 7758 6554 7782 6556
rect 7838 6554 7862 6556
rect 7918 6554 7942 6556
rect 7998 6554 8004 6556
rect 7758 6502 7760 6554
rect 7940 6502 7942 6554
rect 7696 6500 7702 6502
rect 7758 6500 7782 6502
rect 7838 6500 7862 6502
rect 7918 6500 7942 6502
rect 7998 6500 8004 6502
rect 7696 6480 8004 6500
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 7024 5370 7052 5646
rect 7116 5574 7144 6258
rect 7576 5794 7604 6394
rect 7484 5766 7604 5794
rect 8128 5778 8156 6734
rect 8220 6390 8248 6870
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8116 5772 8168 5778
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 5644 4826 5672 5170
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5736 4622 5764 5170
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6010 4924 6318 4944
rect 6010 4922 6016 4924
rect 6072 4922 6096 4924
rect 6152 4922 6176 4924
rect 6232 4922 6256 4924
rect 6312 4922 6318 4924
rect 6072 4870 6074 4922
rect 6254 4870 6256 4922
rect 6010 4868 6016 4870
rect 6072 4868 6096 4870
rect 6152 4868 6176 4870
rect 6232 4868 6256 4870
rect 6312 4868 6318 4870
rect 6010 4848 6318 4868
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 5540 4548 5592 4554
rect 5540 4490 5592 4496
rect 5552 4282 5580 4490
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5736 3738 5764 4558
rect 6380 4078 6408 4558
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 6380 3942 6408 4014
rect 6656 3942 6684 5102
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 7208 4554 7236 4966
rect 7484 4622 7512 5766
rect 8116 5714 8168 5720
rect 8404 5710 8432 6190
rect 8956 5710 8984 7278
rect 9383 7100 9691 7120
rect 9383 7098 9389 7100
rect 9445 7098 9469 7100
rect 9525 7098 9549 7100
rect 9605 7098 9629 7100
rect 9685 7098 9691 7100
rect 9445 7046 9447 7098
rect 9627 7046 9629 7098
rect 9383 7044 9389 7046
rect 9445 7044 9469 7046
rect 9525 7044 9549 7046
rect 9605 7044 9629 7046
rect 9685 7044 9691 7046
rect 9383 7024 9691 7044
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9416 6254 9444 6734
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9036 6248 9088 6254
rect 9036 6190 9088 6196
rect 9404 6248 9456 6254
rect 9404 6190 9456 6196
rect 9048 5778 9076 6190
rect 9383 6012 9691 6032
rect 9383 6010 9389 6012
rect 9445 6010 9469 6012
rect 9525 6010 9549 6012
rect 9605 6010 9629 6012
rect 9685 6010 9691 6012
rect 9445 5958 9447 6010
rect 9627 5958 9629 6010
rect 9383 5956 9389 5958
rect 9445 5956 9469 5958
rect 9525 5956 9549 5958
rect 9605 5956 9629 5958
rect 9685 5956 9691 5958
rect 9383 5936 9691 5956
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 7696 5468 8004 5488
rect 7696 5466 7702 5468
rect 7758 5466 7782 5468
rect 7838 5466 7862 5468
rect 7918 5466 7942 5468
rect 7998 5466 8004 5468
rect 7758 5414 7760 5466
rect 7940 5414 7942 5466
rect 7696 5412 7702 5414
rect 7758 5412 7782 5414
rect 7838 5412 7862 5414
rect 7918 5412 7942 5414
rect 7998 5412 8004 5414
rect 7696 5392 8004 5412
rect 8128 5302 8156 5510
rect 8116 5296 8168 5302
rect 8116 5238 8168 5244
rect 8208 5296 8260 5302
rect 8208 5238 8260 5244
rect 8220 4706 8248 5238
rect 8404 5166 8432 5646
rect 9048 5522 9076 5714
rect 8956 5494 9076 5522
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 8956 5370 8984 5494
rect 8944 5364 8996 5370
rect 8944 5306 8996 5312
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 9383 4924 9691 4944
rect 9383 4922 9389 4924
rect 9445 4922 9469 4924
rect 9525 4922 9549 4924
rect 9605 4922 9629 4924
rect 9685 4922 9691 4924
rect 9445 4870 9447 4922
rect 9627 4870 9629 4922
rect 9383 4868 9389 4870
rect 9445 4868 9469 4870
rect 9525 4868 9549 4870
rect 9605 4868 9629 4870
rect 9685 4868 9691 4870
rect 9383 4848 9691 4868
rect 8036 4690 8248 4706
rect 8036 4684 8260 4690
rect 8036 4678 8208 4684
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7196 4548 7248 4554
rect 7196 4490 7248 4496
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6010 3836 6318 3856
rect 6010 3834 6016 3836
rect 6072 3834 6096 3836
rect 6152 3834 6176 3836
rect 6232 3834 6256 3836
rect 6312 3834 6318 3836
rect 6072 3782 6074 3834
rect 6254 3782 6256 3834
rect 6010 3780 6016 3782
rect 6072 3780 6096 3782
rect 6152 3780 6176 3782
rect 6232 3780 6256 3782
rect 6312 3780 6318 3782
rect 6010 3760 6318 3780
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 6380 3126 6408 3878
rect 6656 3534 6684 3878
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6368 3120 6420 3126
rect 6368 3062 6420 3068
rect 6656 3058 6684 3470
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6010 2748 6318 2768
rect 6010 2746 6016 2748
rect 6072 2746 6096 2748
rect 6152 2746 6176 2748
rect 6232 2746 6256 2748
rect 6312 2746 6318 2748
rect 6072 2694 6074 2746
rect 6254 2694 6256 2746
rect 6010 2692 6016 2694
rect 6072 2692 6096 2694
rect 6152 2692 6176 2694
rect 6232 2692 6256 2694
rect 6312 2692 6318 2694
rect 6010 2672 6318 2692
rect 4252 2576 4304 2582
rect 4252 2518 4304 2524
rect 4160 2508 4212 2514
rect 4160 2450 4212 2456
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 32 800 60 2314
rect 3252 800 3280 2382
rect 4323 2204 4631 2224
rect 4323 2202 4329 2204
rect 4385 2202 4409 2204
rect 4465 2202 4489 2204
rect 4545 2202 4569 2204
rect 4625 2202 4631 2204
rect 4385 2150 4387 2202
rect 4567 2150 4569 2202
rect 4323 2148 4329 2150
rect 4385 2148 4409 2150
rect 4465 2148 4489 2150
rect 4545 2148 4569 2150
rect 4625 2148 4631 2150
rect 4323 2128 4631 2148
rect 6472 800 6500 2790
rect 6656 2514 6684 2994
rect 6932 2514 6960 4422
rect 7208 4078 7236 4490
rect 7484 4282 7512 4558
rect 7696 4380 8004 4400
rect 7696 4378 7702 4380
rect 7758 4378 7782 4380
rect 7838 4378 7862 4380
rect 7918 4378 7942 4380
rect 7998 4378 8004 4380
rect 7758 4326 7760 4378
rect 7940 4326 7942 4378
rect 7696 4324 7702 4326
rect 7758 4324 7782 4326
rect 7838 4324 7862 4326
rect 7918 4324 7942 4326
rect 7998 4324 8004 4326
rect 7696 4304 8004 4324
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 8036 3534 8064 4678
rect 8208 4626 8260 4632
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 8208 4548 8260 4554
rect 8208 4490 8260 4496
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 7696 3292 8004 3312
rect 7696 3290 7702 3292
rect 7758 3290 7782 3292
rect 7838 3290 7862 3292
rect 7918 3290 7942 3292
rect 7998 3290 8004 3292
rect 7758 3238 7760 3290
rect 7940 3238 7942 3290
rect 7696 3236 7702 3238
rect 7758 3236 7782 3238
rect 7838 3236 7862 3238
rect 7918 3236 7942 3238
rect 7998 3236 8004 3238
rect 7696 3216 8004 3236
rect 8036 3126 8064 3470
rect 8024 3120 8076 3126
rect 8024 3062 8076 3068
rect 6644 2508 6696 2514
rect 6644 2450 6696 2456
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 8036 2446 8064 3062
rect 8220 2650 8248 4490
rect 9324 4214 9352 4626
rect 9312 4208 9364 4214
rect 9312 4150 9364 4156
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 9048 3194 9076 4014
rect 9383 3836 9691 3856
rect 9383 3834 9389 3836
rect 9445 3834 9469 3836
rect 9525 3834 9549 3836
rect 9605 3834 9629 3836
rect 9685 3834 9691 3836
rect 9445 3782 9447 3834
rect 9627 3782 9629 3834
rect 9383 3780 9389 3782
rect 9445 3780 9469 3782
rect 9525 3780 9549 3782
rect 9605 3780 9629 3782
rect 9685 3780 9691 3782
rect 9383 3760 9691 3780
rect 9784 3670 9812 5510
rect 9772 3664 9824 3670
rect 9772 3606 9824 3612
rect 9876 3602 9904 6598
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 9968 3534 9996 10542
rect 10060 10266 10088 11086
rect 10152 10810 10180 11154
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 10244 8906 10272 11086
rect 10428 10985 10456 11222
rect 10414 10976 10470 10985
rect 10414 10911 10470 10920
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10336 10062 10364 10406
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10232 8900 10284 8906
rect 10232 8842 10284 8848
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 10428 7585 10456 7686
rect 10414 7576 10470 7585
rect 10414 7511 10470 7520
rect 10232 7336 10284 7342
rect 10232 7278 10284 7284
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10140 6724 10192 6730
rect 10140 6666 10192 6672
rect 10152 5302 10180 6666
rect 10244 6458 10272 7278
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10140 5296 10192 5302
rect 10140 5238 10192 5244
rect 10324 5296 10376 5302
rect 10324 5238 10376 5244
rect 10336 4282 10364 5238
rect 10520 5234 10548 7278
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10324 4276 10376 4282
rect 10324 4218 10376 4224
rect 10520 4185 10548 4558
rect 10506 4176 10562 4185
rect 10506 4111 10562 4120
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 9383 2748 9691 2768
rect 9383 2746 9389 2748
rect 9445 2746 9469 2748
rect 9525 2746 9549 2748
rect 9605 2746 9629 2748
rect 9685 2746 9691 2748
rect 9445 2694 9447 2746
rect 9627 2694 9629 2746
rect 9383 2692 9389 2694
rect 9445 2692 9469 2694
rect 9525 2692 9549 2694
rect 9605 2692 9629 2694
rect 9685 2692 9691 2694
rect 9383 2672 9691 2692
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 9968 2446 9996 3470
rect 8024 2440 8076 2446
rect 8024 2382 8076 2388
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 10416 2304 10468 2310
rect 10416 2246 10468 2252
rect 7696 2204 8004 2224
rect 7696 2202 7702 2204
rect 7758 2202 7782 2204
rect 7838 2202 7862 2204
rect 7918 2202 7942 2204
rect 7998 2202 8004 2204
rect 7758 2150 7760 2202
rect 7940 2150 7942 2202
rect 7696 2148 7702 2150
rect 7758 2148 7782 2150
rect 7838 2148 7862 2150
rect 7918 2148 7942 2150
rect 7998 2148 8004 2150
rect 7696 2128 8004 2148
rect 9692 800 9720 2246
rect 18 0 74 800
rect 3238 0 3294 800
rect 6458 0 6514 800
rect 9678 0 9734 800
rect 10428 785 10456 2246
rect 10414 776 10470 785
rect 10414 711 10470 720
<< via2 >>
rect 1490 13640 1546 13696
rect 4329 11994 4385 11996
rect 4409 11994 4465 11996
rect 4489 11994 4545 11996
rect 4569 11994 4625 11996
rect 4329 11942 4375 11994
rect 4375 11942 4385 11994
rect 4409 11942 4439 11994
rect 4439 11942 4451 11994
rect 4451 11942 4465 11994
rect 4489 11942 4503 11994
rect 4503 11942 4515 11994
rect 4515 11942 4545 11994
rect 4569 11942 4579 11994
rect 4579 11942 4625 11994
rect 4329 11940 4385 11942
rect 4409 11940 4465 11942
rect 4489 11940 4545 11942
rect 4569 11940 4625 11942
rect 7702 11994 7758 11996
rect 7782 11994 7838 11996
rect 7862 11994 7918 11996
rect 7942 11994 7998 11996
rect 7702 11942 7748 11994
rect 7748 11942 7758 11994
rect 7782 11942 7812 11994
rect 7812 11942 7824 11994
rect 7824 11942 7838 11994
rect 7862 11942 7876 11994
rect 7876 11942 7888 11994
rect 7888 11942 7918 11994
rect 7942 11942 7952 11994
rect 7952 11942 7998 11994
rect 7702 11940 7758 11942
rect 7782 11940 7838 11942
rect 7862 11940 7918 11942
rect 7942 11940 7998 11942
rect 1490 10260 1546 10296
rect 1490 10240 1492 10260
rect 1492 10240 1544 10260
rect 1544 10240 1546 10260
rect 1490 6876 1492 6896
rect 1492 6876 1544 6896
rect 1544 6876 1546 6896
rect 1490 6840 1546 6876
rect 2642 11450 2698 11452
rect 2722 11450 2778 11452
rect 2802 11450 2858 11452
rect 2882 11450 2938 11452
rect 2642 11398 2688 11450
rect 2688 11398 2698 11450
rect 2722 11398 2752 11450
rect 2752 11398 2764 11450
rect 2764 11398 2778 11450
rect 2802 11398 2816 11450
rect 2816 11398 2828 11450
rect 2828 11398 2858 11450
rect 2882 11398 2892 11450
rect 2892 11398 2938 11450
rect 2642 11396 2698 11398
rect 2722 11396 2778 11398
rect 2802 11396 2858 11398
rect 2882 11396 2938 11398
rect 2642 10362 2698 10364
rect 2722 10362 2778 10364
rect 2802 10362 2858 10364
rect 2882 10362 2938 10364
rect 2642 10310 2688 10362
rect 2688 10310 2698 10362
rect 2722 10310 2752 10362
rect 2752 10310 2764 10362
rect 2764 10310 2778 10362
rect 2802 10310 2816 10362
rect 2816 10310 2828 10362
rect 2828 10310 2858 10362
rect 2882 10310 2892 10362
rect 2892 10310 2938 10362
rect 2642 10308 2698 10310
rect 2722 10308 2778 10310
rect 2802 10308 2858 10310
rect 2882 10308 2938 10310
rect 4329 10906 4385 10908
rect 4409 10906 4465 10908
rect 4489 10906 4545 10908
rect 4569 10906 4625 10908
rect 4329 10854 4375 10906
rect 4375 10854 4385 10906
rect 4409 10854 4439 10906
rect 4439 10854 4451 10906
rect 4451 10854 4465 10906
rect 4489 10854 4503 10906
rect 4503 10854 4515 10906
rect 4515 10854 4545 10906
rect 4569 10854 4579 10906
rect 4579 10854 4625 10906
rect 4329 10852 4385 10854
rect 4409 10852 4465 10854
rect 4489 10852 4545 10854
rect 4569 10852 4625 10854
rect 4329 9818 4385 9820
rect 4409 9818 4465 9820
rect 4489 9818 4545 9820
rect 4569 9818 4625 9820
rect 4329 9766 4375 9818
rect 4375 9766 4385 9818
rect 4409 9766 4439 9818
rect 4439 9766 4451 9818
rect 4451 9766 4465 9818
rect 4489 9766 4503 9818
rect 4503 9766 4515 9818
rect 4515 9766 4545 9818
rect 4569 9766 4579 9818
rect 4579 9766 4625 9818
rect 4329 9764 4385 9766
rect 4409 9764 4465 9766
rect 4489 9764 4545 9766
rect 4569 9764 4625 9766
rect 2642 9274 2698 9276
rect 2722 9274 2778 9276
rect 2802 9274 2858 9276
rect 2882 9274 2938 9276
rect 2642 9222 2688 9274
rect 2688 9222 2698 9274
rect 2722 9222 2752 9274
rect 2752 9222 2764 9274
rect 2764 9222 2778 9274
rect 2802 9222 2816 9274
rect 2816 9222 2828 9274
rect 2828 9222 2858 9274
rect 2882 9222 2892 9274
rect 2892 9222 2938 9274
rect 2642 9220 2698 9222
rect 2722 9220 2778 9222
rect 2802 9220 2858 9222
rect 2882 9220 2938 9222
rect 2642 8186 2698 8188
rect 2722 8186 2778 8188
rect 2802 8186 2858 8188
rect 2882 8186 2938 8188
rect 2642 8134 2688 8186
rect 2688 8134 2698 8186
rect 2722 8134 2752 8186
rect 2752 8134 2764 8186
rect 2764 8134 2778 8186
rect 2802 8134 2816 8186
rect 2816 8134 2828 8186
rect 2828 8134 2858 8186
rect 2882 8134 2892 8186
rect 2892 8134 2938 8186
rect 2642 8132 2698 8134
rect 2722 8132 2778 8134
rect 2802 8132 2858 8134
rect 2882 8132 2938 8134
rect 2642 7098 2698 7100
rect 2722 7098 2778 7100
rect 2802 7098 2858 7100
rect 2882 7098 2938 7100
rect 2642 7046 2688 7098
rect 2688 7046 2698 7098
rect 2722 7046 2752 7098
rect 2752 7046 2764 7098
rect 2764 7046 2778 7098
rect 2802 7046 2816 7098
rect 2816 7046 2828 7098
rect 2828 7046 2858 7098
rect 2882 7046 2892 7098
rect 2892 7046 2938 7098
rect 2642 7044 2698 7046
rect 2722 7044 2778 7046
rect 2802 7044 2858 7046
rect 2882 7044 2938 7046
rect 4329 8730 4385 8732
rect 4409 8730 4465 8732
rect 4489 8730 4545 8732
rect 4569 8730 4625 8732
rect 4329 8678 4375 8730
rect 4375 8678 4385 8730
rect 4409 8678 4439 8730
rect 4439 8678 4451 8730
rect 4451 8678 4465 8730
rect 4489 8678 4503 8730
rect 4503 8678 4515 8730
rect 4515 8678 4545 8730
rect 4569 8678 4579 8730
rect 4579 8678 4625 8730
rect 4329 8676 4385 8678
rect 4409 8676 4465 8678
rect 4489 8676 4545 8678
rect 4569 8676 4625 8678
rect 4329 7642 4385 7644
rect 4409 7642 4465 7644
rect 4489 7642 4545 7644
rect 4569 7642 4625 7644
rect 4329 7590 4375 7642
rect 4375 7590 4385 7642
rect 4409 7590 4439 7642
rect 4439 7590 4451 7642
rect 4451 7590 4465 7642
rect 4489 7590 4503 7642
rect 4503 7590 4515 7642
rect 4515 7590 4545 7642
rect 4569 7590 4579 7642
rect 4579 7590 4625 7642
rect 4329 7588 4385 7590
rect 4409 7588 4465 7590
rect 4489 7588 4545 7590
rect 4569 7588 4625 7590
rect 4329 6554 4385 6556
rect 4409 6554 4465 6556
rect 4489 6554 4545 6556
rect 4569 6554 4625 6556
rect 4329 6502 4375 6554
rect 4375 6502 4385 6554
rect 4409 6502 4439 6554
rect 4439 6502 4451 6554
rect 4451 6502 4465 6554
rect 4489 6502 4503 6554
rect 4503 6502 4515 6554
rect 4515 6502 4545 6554
rect 4569 6502 4579 6554
rect 4579 6502 4625 6554
rect 4329 6500 4385 6502
rect 4409 6500 4465 6502
rect 4489 6500 4545 6502
rect 4569 6500 4625 6502
rect 2642 6010 2698 6012
rect 2722 6010 2778 6012
rect 2802 6010 2858 6012
rect 2882 6010 2938 6012
rect 2642 5958 2688 6010
rect 2688 5958 2698 6010
rect 2722 5958 2752 6010
rect 2752 5958 2764 6010
rect 2764 5958 2778 6010
rect 2802 5958 2816 6010
rect 2816 5958 2828 6010
rect 2828 5958 2858 6010
rect 2882 5958 2892 6010
rect 2892 5958 2938 6010
rect 2642 5956 2698 5958
rect 2722 5956 2778 5958
rect 2802 5956 2858 5958
rect 2882 5956 2938 5958
rect 2642 4922 2698 4924
rect 2722 4922 2778 4924
rect 2802 4922 2858 4924
rect 2882 4922 2938 4924
rect 2642 4870 2688 4922
rect 2688 4870 2698 4922
rect 2722 4870 2752 4922
rect 2752 4870 2764 4922
rect 2764 4870 2778 4922
rect 2802 4870 2816 4922
rect 2816 4870 2828 4922
rect 2828 4870 2858 4922
rect 2882 4870 2892 4922
rect 2892 4870 2938 4922
rect 2642 4868 2698 4870
rect 2722 4868 2778 4870
rect 2802 4868 2858 4870
rect 2882 4868 2938 4870
rect 1490 3440 1546 3496
rect 4329 5466 4385 5468
rect 4409 5466 4465 5468
rect 4489 5466 4545 5468
rect 4569 5466 4625 5468
rect 4329 5414 4375 5466
rect 4375 5414 4385 5466
rect 4409 5414 4439 5466
rect 4439 5414 4451 5466
rect 4451 5414 4465 5466
rect 4489 5414 4503 5466
rect 4503 5414 4515 5466
rect 4515 5414 4545 5466
rect 4569 5414 4579 5466
rect 4579 5414 4625 5466
rect 4329 5412 4385 5414
rect 4409 5412 4465 5414
rect 4489 5412 4545 5414
rect 4569 5412 4625 5414
rect 2642 3834 2698 3836
rect 2722 3834 2778 3836
rect 2802 3834 2858 3836
rect 2882 3834 2938 3836
rect 2642 3782 2688 3834
rect 2688 3782 2698 3834
rect 2722 3782 2752 3834
rect 2752 3782 2764 3834
rect 2764 3782 2778 3834
rect 2802 3782 2816 3834
rect 2816 3782 2828 3834
rect 2828 3782 2858 3834
rect 2882 3782 2892 3834
rect 2892 3782 2938 3834
rect 2642 3780 2698 3782
rect 2722 3780 2778 3782
rect 2802 3780 2858 3782
rect 2882 3780 2938 3782
rect 4329 4378 4385 4380
rect 4409 4378 4465 4380
rect 4489 4378 4545 4380
rect 4569 4378 4625 4380
rect 4329 4326 4375 4378
rect 4375 4326 4385 4378
rect 4409 4326 4439 4378
rect 4439 4326 4451 4378
rect 4451 4326 4465 4378
rect 4489 4326 4503 4378
rect 4503 4326 4515 4378
rect 4515 4326 4545 4378
rect 4569 4326 4579 4378
rect 4579 4326 4625 4378
rect 4329 4324 4385 4326
rect 4409 4324 4465 4326
rect 4489 4324 4545 4326
rect 4569 4324 4625 4326
rect 2642 2746 2698 2748
rect 2722 2746 2778 2748
rect 2802 2746 2858 2748
rect 2882 2746 2938 2748
rect 2642 2694 2688 2746
rect 2688 2694 2698 2746
rect 2722 2694 2752 2746
rect 2752 2694 2764 2746
rect 2764 2694 2778 2746
rect 2802 2694 2816 2746
rect 2816 2694 2828 2746
rect 2828 2694 2858 2746
rect 2882 2694 2892 2746
rect 2892 2694 2938 2746
rect 2642 2692 2698 2694
rect 2722 2692 2778 2694
rect 2802 2692 2858 2694
rect 2882 2692 2938 2694
rect 4329 3290 4385 3292
rect 4409 3290 4465 3292
rect 4489 3290 4545 3292
rect 4569 3290 4625 3292
rect 4329 3238 4375 3290
rect 4375 3238 4385 3290
rect 4409 3238 4439 3290
rect 4439 3238 4451 3290
rect 4451 3238 4465 3290
rect 4489 3238 4503 3290
rect 4503 3238 4515 3290
rect 4515 3238 4545 3290
rect 4569 3238 4579 3290
rect 4579 3238 4625 3290
rect 4329 3236 4385 3238
rect 4409 3236 4465 3238
rect 4489 3236 4545 3238
rect 4569 3236 4625 3238
rect 6016 11450 6072 11452
rect 6096 11450 6152 11452
rect 6176 11450 6232 11452
rect 6256 11450 6312 11452
rect 6016 11398 6062 11450
rect 6062 11398 6072 11450
rect 6096 11398 6126 11450
rect 6126 11398 6138 11450
rect 6138 11398 6152 11450
rect 6176 11398 6190 11450
rect 6190 11398 6202 11450
rect 6202 11398 6232 11450
rect 6256 11398 6266 11450
rect 6266 11398 6312 11450
rect 6016 11396 6072 11398
rect 6096 11396 6152 11398
rect 6176 11396 6232 11398
rect 6256 11396 6312 11398
rect 7702 10906 7758 10908
rect 7782 10906 7838 10908
rect 7862 10906 7918 10908
rect 7942 10906 7998 10908
rect 7702 10854 7748 10906
rect 7748 10854 7758 10906
rect 7782 10854 7812 10906
rect 7812 10854 7824 10906
rect 7824 10854 7838 10906
rect 7862 10854 7876 10906
rect 7876 10854 7888 10906
rect 7888 10854 7918 10906
rect 7942 10854 7952 10906
rect 7952 10854 7998 10906
rect 7702 10852 7758 10854
rect 7782 10852 7838 10854
rect 7862 10852 7918 10854
rect 7942 10852 7998 10854
rect 6016 10362 6072 10364
rect 6096 10362 6152 10364
rect 6176 10362 6232 10364
rect 6256 10362 6312 10364
rect 6016 10310 6062 10362
rect 6062 10310 6072 10362
rect 6096 10310 6126 10362
rect 6126 10310 6138 10362
rect 6138 10310 6152 10362
rect 6176 10310 6190 10362
rect 6190 10310 6202 10362
rect 6202 10310 6232 10362
rect 6256 10310 6266 10362
rect 6266 10310 6312 10362
rect 6016 10308 6072 10310
rect 6096 10308 6152 10310
rect 6176 10308 6232 10310
rect 6256 10308 6312 10310
rect 6016 9274 6072 9276
rect 6096 9274 6152 9276
rect 6176 9274 6232 9276
rect 6256 9274 6312 9276
rect 6016 9222 6062 9274
rect 6062 9222 6072 9274
rect 6096 9222 6126 9274
rect 6126 9222 6138 9274
rect 6138 9222 6152 9274
rect 6176 9222 6190 9274
rect 6190 9222 6202 9274
rect 6202 9222 6232 9274
rect 6256 9222 6266 9274
rect 6266 9222 6312 9274
rect 6016 9220 6072 9222
rect 6096 9220 6152 9222
rect 6176 9220 6232 9222
rect 6256 9220 6312 9222
rect 6016 8186 6072 8188
rect 6096 8186 6152 8188
rect 6176 8186 6232 8188
rect 6256 8186 6312 8188
rect 6016 8134 6062 8186
rect 6062 8134 6072 8186
rect 6096 8134 6126 8186
rect 6126 8134 6138 8186
rect 6138 8134 6152 8186
rect 6176 8134 6190 8186
rect 6190 8134 6202 8186
rect 6202 8134 6232 8186
rect 6256 8134 6266 8186
rect 6266 8134 6312 8186
rect 6016 8132 6072 8134
rect 6096 8132 6152 8134
rect 6176 8132 6232 8134
rect 6256 8132 6312 8134
rect 7702 9818 7758 9820
rect 7782 9818 7838 9820
rect 7862 9818 7918 9820
rect 7942 9818 7998 9820
rect 7702 9766 7748 9818
rect 7748 9766 7758 9818
rect 7782 9766 7812 9818
rect 7812 9766 7824 9818
rect 7824 9766 7838 9818
rect 7862 9766 7876 9818
rect 7876 9766 7888 9818
rect 7888 9766 7918 9818
rect 7942 9766 7952 9818
rect 7952 9766 7998 9818
rect 7702 9764 7758 9766
rect 7782 9764 7838 9766
rect 7862 9764 7918 9766
rect 7942 9764 7998 9766
rect 7702 8730 7758 8732
rect 7782 8730 7838 8732
rect 7862 8730 7918 8732
rect 7942 8730 7998 8732
rect 7702 8678 7748 8730
rect 7748 8678 7758 8730
rect 7782 8678 7812 8730
rect 7812 8678 7824 8730
rect 7824 8678 7838 8730
rect 7862 8678 7876 8730
rect 7876 8678 7888 8730
rect 7888 8678 7918 8730
rect 7942 8678 7952 8730
rect 7952 8678 7998 8730
rect 7702 8676 7758 8678
rect 7782 8676 7838 8678
rect 7862 8676 7918 8678
rect 7942 8676 7998 8678
rect 9389 11450 9445 11452
rect 9469 11450 9525 11452
rect 9549 11450 9605 11452
rect 9629 11450 9685 11452
rect 9389 11398 9435 11450
rect 9435 11398 9445 11450
rect 9469 11398 9499 11450
rect 9499 11398 9511 11450
rect 9511 11398 9525 11450
rect 9549 11398 9563 11450
rect 9563 11398 9575 11450
rect 9575 11398 9605 11450
rect 9629 11398 9639 11450
rect 9639 11398 9685 11450
rect 9389 11396 9445 11398
rect 9469 11396 9525 11398
rect 9549 11396 9605 11398
rect 9629 11396 9685 11398
rect 9389 10362 9445 10364
rect 9469 10362 9525 10364
rect 9549 10362 9605 10364
rect 9629 10362 9685 10364
rect 9389 10310 9435 10362
rect 9435 10310 9445 10362
rect 9469 10310 9499 10362
rect 9499 10310 9511 10362
rect 9511 10310 9525 10362
rect 9549 10310 9563 10362
rect 9563 10310 9575 10362
rect 9575 10310 9605 10362
rect 9629 10310 9639 10362
rect 9639 10310 9685 10362
rect 9389 10308 9445 10310
rect 9469 10308 9525 10310
rect 9549 10308 9605 10310
rect 9629 10308 9685 10310
rect 6016 7098 6072 7100
rect 6096 7098 6152 7100
rect 6176 7098 6232 7100
rect 6256 7098 6312 7100
rect 6016 7046 6062 7098
rect 6062 7046 6072 7098
rect 6096 7046 6126 7098
rect 6126 7046 6138 7098
rect 6138 7046 6152 7098
rect 6176 7046 6190 7098
rect 6190 7046 6202 7098
rect 6202 7046 6232 7098
rect 6256 7046 6266 7098
rect 6266 7046 6312 7098
rect 6016 7044 6072 7046
rect 6096 7044 6152 7046
rect 6176 7044 6232 7046
rect 6256 7044 6312 7046
rect 6016 6010 6072 6012
rect 6096 6010 6152 6012
rect 6176 6010 6232 6012
rect 6256 6010 6312 6012
rect 6016 5958 6062 6010
rect 6062 5958 6072 6010
rect 6096 5958 6126 6010
rect 6126 5958 6138 6010
rect 6138 5958 6152 6010
rect 6176 5958 6190 6010
rect 6190 5958 6202 6010
rect 6202 5958 6232 6010
rect 6256 5958 6266 6010
rect 6266 5958 6312 6010
rect 6016 5956 6072 5958
rect 6096 5956 6152 5958
rect 6176 5956 6232 5958
rect 6256 5956 6312 5958
rect 7702 7642 7758 7644
rect 7782 7642 7838 7644
rect 7862 7642 7918 7644
rect 7942 7642 7998 7644
rect 7702 7590 7748 7642
rect 7748 7590 7758 7642
rect 7782 7590 7812 7642
rect 7812 7590 7824 7642
rect 7824 7590 7838 7642
rect 7862 7590 7876 7642
rect 7876 7590 7888 7642
rect 7888 7590 7918 7642
rect 7942 7590 7952 7642
rect 7952 7590 7998 7642
rect 7702 7588 7758 7590
rect 7782 7588 7838 7590
rect 7862 7588 7918 7590
rect 7942 7588 7998 7590
rect 9389 9274 9445 9276
rect 9469 9274 9525 9276
rect 9549 9274 9605 9276
rect 9629 9274 9685 9276
rect 9389 9222 9435 9274
rect 9435 9222 9445 9274
rect 9469 9222 9499 9274
rect 9499 9222 9511 9274
rect 9511 9222 9525 9274
rect 9549 9222 9563 9274
rect 9563 9222 9575 9274
rect 9575 9222 9605 9274
rect 9629 9222 9639 9274
rect 9639 9222 9685 9274
rect 9389 9220 9445 9222
rect 9469 9220 9525 9222
rect 9549 9220 9605 9222
rect 9629 9220 9685 9222
rect 9389 8186 9445 8188
rect 9469 8186 9525 8188
rect 9549 8186 9605 8188
rect 9629 8186 9685 8188
rect 9389 8134 9435 8186
rect 9435 8134 9445 8186
rect 9469 8134 9499 8186
rect 9499 8134 9511 8186
rect 9511 8134 9525 8186
rect 9549 8134 9563 8186
rect 9563 8134 9575 8186
rect 9575 8134 9605 8186
rect 9629 8134 9639 8186
rect 9639 8134 9685 8186
rect 9389 8132 9445 8134
rect 9469 8132 9525 8134
rect 9549 8132 9605 8134
rect 9629 8132 9685 8134
rect 7702 6554 7758 6556
rect 7782 6554 7838 6556
rect 7862 6554 7918 6556
rect 7942 6554 7998 6556
rect 7702 6502 7748 6554
rect 7748 6502 7758 6554
rect 7782 6502 7812 6554
rect 7812 6502 7824 6554
rect 7824 6502 7838 6554
rect 7862 6502 7876 6554
rect 7876 6502 7888 6554
rect 7888 6502 7918 6554
rect 7942 6502 7952 6554
rect 7952 6502 7998 6554
rect 7702 6500 7758 6502
rect 7782 6500 7838 6502
rect 7862 6500 7918 6502
rect 7942 6500 7998 6502
rect 6016 4922 6072 4924
rect 6096 4922 6152 4924
rect 6176 4922 6232 4924
rect 6256 4922 6312 4924
rect 6016 4870 6062 4922
rect 6062 4870 6072 4922
rect 6096 4870 6126 4922
rect 6126 4870 6138 4922
rect 6138 4870 6152 4922
rect 6176 4870 6190 4922
rect 6190 4870 6202 4922
rect 6202 4870 6232 4922
rect 6256 4870 6266 4922
rect 6266 4870 6312 4922
rect 6016 4868 6072 4870
rect 6096 4868 6152 4870
rect 6176 4868 6232 4870
rect 6256 4868 6312 4870
rect 9389 7098 9445 7100
rect 9469 7098 9525 7100
rect 9549 7098 9605 7100
rect 9629 7098 9685 7100
rect 9389 7046 9435 7098
rect 9435 7046 9445 7098
rect 9469 7046 9499 7098
rect 9499 7046 9511 7098
rect 9511 7046 9525 7098
rect 9549 7046 9563 7098
rect 9563 7046 9575 7098
rect 9575 7046 9605 7098
rect 9629 7046 9639 7098
rect 9639 7046 9685 7098
rect 9389 7044 9445 7046
rect 9469 7044 9525 7046
rect 9549 7044 9605 7046
rect 9629 7044 9685 7046
rect 9389 6010 9445 6012
rect 9469 6010 9525 6012
rect 9549 6010 9605 6012
rect 9629 6010 9685 6012
rect 9389 5958 9435 6010
rect 9435 5958 9445 6010
rect 9469 5958 9499 6010
rect 9499 5958 9511 6010
rect 9511 5958 9525 6010
rect 9549 5958 9563 6010
rect 9563 5958 9575 6010
rect 9575 5958 9605 6010
rect 9629 5958 9639 6010
rect 9639 5958 9685 6010
rect 9389 5956 9445 5958
rect 9469 5956 9525 5958
rect 9549 5956 9605 5958
rect 9629 5956 9685 5958
rect 7702 5466 7758 5468
rect 7782 5466 7838 5468
rect 7862 5466 7918 5468
rect 7942 5466 7998 5468
rect 7702 5414 7748 5466
rect 7748 5414 7758 5466
rect 7782 5414 7812 5466
rect 7812 5414 7824 5466
rect 7824 5414 7838 5466
rect 7862 5414 7876 5466
rect 7876 5414 7888 5466
rect 7888 5414 7918 5466
rect 7942 5414 7952 5466
rect 7952 5414 7998 5466
rect 7702 5412 7758 5414
rect 7782 5412 7838 5414
rect 7862 5412 7918 5414
rect 7942 5412 7998 5414
rect 9389 4922 9445 4924
rect 9469 4922 9525 4924
rect 9549 4922 9605 4924
rect 9629 4922 9685 4924
rect 9389 4870 9435 4922
rect 9435 4870 9445 4922
rect 9469 4870 9499 4922
rect 9499 4870 9511 4922
rect 9511 4870 9525 4922
rect 9549 4870 9563 4922
rect 9563 4870 9575 4922
rect 9575 4870 9605 4922
rect 9629 4870 9639 4922
rect 9639 4870 9685 4922
rect 9389 4868 9445 4870
rect 9469 4868 9525 4870
rect 9549 4868 9605 4870
rect 9629 4868 9685 4870
rect 6016 3834 6072 3836
rect 6096 3834 6152 3836
rect 6176 3834 6232 3836
rect 6256 3834 6312 3836
rect 6016 3782 6062 3834
rect 6062 3782 6072 3834
rect 6096 3782 6126 3834
rect 6126 3782 6138 3834
rect 6138 3782 6152 3834
rect 6176 3782 6190 3834
rect 6190 3782 6202 3834
rect 6202 3782 6232 3834
rect 6256 3782 6266 3834
rect 6266 3782 6312 3834
rect 6016 3780 6072 3782
rect 6096 3780 6152 3782
rect 6176 3780 6232 3782
rect 6256 3780 6312 3782
rect 6016 2746 6072 2748
rect 6096 2746 6152 2748
rect 6176 2746 6232 2748
rect 6256 2746 6312 2748
rect 6016 2694 6062 2746
rect 6062 2694 6072 2746
rect 6096 2694 6126 2746
rect 6126 2694 6138 2746
rect 6138 2694 6152 2746
rect 6176 2694 6190 2746
rect 6190 2694 6202 2746
rect 6202 2694 6232 2746
rect 6256 2694 6266 2746
rect 6266 2694 6312 2746
rect 6016 2692 6072 2694
rect 6096 2692 6152 2694
rect 6176 2692 6232 2694
rect 6256 2692 6312 2694
rect 4329 2202 4385 2204
rect 4409 2202 4465 2204
rect 4489 2202 4545 2204
rect 4569 2202 4625 2204
rect 4329 2150 4375 2202
rect 4375 2150 4385 2202
rect 4409 2150 4439 2202
rect 4439 2150 4451 2202
rect 4451 2150 4465 2202
rect 4489 2150 4503 2202
rect 4503 2150 4515 2202
rect 4515 2150 4545 2202
rect 4569 2150 4579 2202
rect 4579 2150 4625 2202
rect 4329 2148 4385 2150
rect 4409 2148 4465 2150
rect 4489 2148 4545 2150
rect 4569 2148 4625 2150
rect 7702 4378 7758 4380
rect 7782 4378 7838 4380
rect 7862 4378 7918 4380
rect 7942 4378 7998 4380
rect 7702 4326 7748 4378
rect 7748 4326 7758 4378
rect 7782 4326 7812 4378
rect 7812 4326 7824 4378
rect 7824 4326 7838 4378
rect 7862 4326 7876 4378
rect 7876 4326 7888 4378
rect 7888 4326 7918 4378
rect 7942 4326 7952 4378
rect 7952 4326 7998 4378
rect 7702 4324 7758 4326
rect 7782 4324 7838 4326
rect 7862 4324 7918 4326
rect 7942 4324 7998 4326
rect 7702 3290 7758 3292
rect 7782 3290 7838 3292
rect 7862 3290 7918 3292
rect 7942 3290 7998 3292
rect 7702 3238 7748 3290
rect 7748 3238 7758 3290
rect 7782 3238 7812 3290
rect 7812 3238 7824 3290
rect 7824 3238 7838 3290
rect 7862 3238 7876 3290
rect 7876 3238 7888 3290
rect 7888 3238 7918 3290
rect 7942 3238 7952 3290
rect 7952 3238 7998 3290
rect 7702 3236 7758 3238
rect 7782 3236 7838 3238
rect 7862 3236 7918 3238
rect 7942 3236 7998 3238
rect 9389 3834 9445 3836
rect 9469 3834 9525 3836
rect 9549 3834 9605 3836
rect 9629 3834 9685 3836
rect 9389 3782 9435 3834
rect 9435 3782 9445 3834
rect 9469 3782 9499 3834
rect 9499 3782 9511 3834
rect 9511 3782 9525 3834
rect 9549 3782 9563 3834
rect 9563 3782 9575 3834
rect 9575 3782 9605 3834
rect 9629 3782 9639 3834
rect 9639 3782 9685 3834
rect 9389 3780 9445 3782
rect 9469 3780 9525 3782
rect 9549 3780 9605 3782
rect 9629 3780 9685 3782
rect 10414 10920 10470 10976
rect 10414 7520 10470 7576
rect 10506 4120 10562 4176
rect 9389 2746 9445 2748
rect 9469 2746 9525 2748
rect 9549 2746 9605 2748
rect 9629 2746 9685 2748
rect 9389 2694 9435 2746
rect 9435 2694 9445 2746
rect 9469 2694 9499 2746
rect 9499 2694 9511 2746
rect 9511 2694 9525 2746
rect 9549 2694 9563 2746
rect 9563 2694 9575 2746
rect 9575 2694 9605 2746
rect 9629 2694 9639 2746
rect 9639 2694 9685 2746
rect 9389 2692 9445 2694
rect 9469 2692 9525 2694
rect 9549 2692 9605 2694
rect 9629 2692 9685 2694
rect 7702 2202 7758 2204
rect 7782 2202 7838 2204
rect 7862 2202 7918 2204
rect 7942 2202 7998 2204
rect 7702 2150 7748 2202
rect 7748 2150 7758 2202
rect 7782 2150 7812 2202
rect 7812 2150 7824 2202
rect 7824 2150 7838 2202
rect 7862 2150 7876 2202
rect 7876 2150 7888 2202
rect 7888 2150 7918 2202
rect 7942 2150 7952 2202
rect 7952 2150 7998 2202
rect 7702 2148 7758 2150
rect 7782 2148 7838 2150
rect 7862 2148 7918 2150
rect 7942 2148 7998 2150
rect 10414 720 10470 776
<< metal3 >>
rect 0 13698 800 13728
rect 1485 13698 1551 13701
rect 0 13696 1551 13698
rect 0 13640 1490 13696
rect 1546 13640 1551 13696
rect 0 13638 1551 13640
rect 0 13608 800 13638
rect 1485 13635 1551 13638
rect 4317 12000 4637 12001
rect 4317 11936 4325 12000
rect 4389 11936 4405 12000
rect 4469 11936 4485 12000
rect 4549 11936 4565 12000
rect 4629 11936 4637 12000
rect 4317 11935 4637 11936
rect 7690 12000 8010 12001
rect 7690 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7938 12000
rect 8002 11936 8010 12000
rect 7690 11935 8010 11936
rect 2630 11456 2950 11457
rect 2630 11392 2638 11456
rect 2702 11392 2718 11456
rect 2782 11392 2798 11456
rect 2862 11392 2878 11456
rect 2942 11392 2950 11456
rect 2630 11391 2950 11392
rect 6004 11456 6324 11457
rect 6004 11392 6012 11456
rect 6076 11392 6092 11456
rect 6156 11392 6172 11456
rect 6236 11392 6252 11456
rect 6316 11392 6324 11456
rect 6004 11391 6324 11392
rect 9377 11456 9697 11457
rect 9377 11392 9385 11456
rect 9449 11392 9465 11456
rect 9529 11392 9545 11456
rect 9609 11392 9625 11456
rect 9689 11392 9697 11456
rect 9377 11391 9697 11392
rect 10409 10978 10475 10981
rect 11529 10978 12329 11008
rect 10409 10976 12329 10978
rect 10409 10920 10414 10976
rect 10470 10920 12329 10976
rect 10409 10918 12329 10920
rect 10409 10915 10475 10918
rect 4317 10912 4637 10913
rect 4317 10848 4325 10912
rect 4389 10848 4405 10912
rect 4469 10848 4485 10912
rect 4549 10848 4565 10912
rect 4629 10848 4637 10912
rect 4317 10847 4637 10848
rect 7690 10912 8010 10913
rect 7690 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7938 10912
rect 8002 10848 8010 10912
rect 11529 10888 12329 10918
rect 7690 10847 8010 10848
rect 2630 10368 2950 10369
rect 0 10298 800 10328
rect 2630 10304 2638 10368
rect 2702 10304 2718 10368
rect 2782 10304 2798 10368
rect 2862 10304 2878 10368
rect 2942 10304 2950 10368
rect 2630 10303 2950 10304
rect 6004 10368 6324 10369
rect 6004 10304 6012 10368
rect 6076 10304 6092 10368
rect 6156 10304 6172 10368
rect 6236 10304 6252 10368
rect 6316 10304 6324 10368
rect 6004 10303 6324 10304
rect 9377 10368 9697 10369
rect 9377 10304 9385 10368
rect 9449 10304 9465 10368
rect 9529 10304 9545 10368
rect 9609 10304 9625 10368
rect 9689 10304 9697 10368
rect 9377 10303 9697 10304
rect 1485 10298 1551 10301
rect 0 10296 1551 10298
rect 0 10240 1490 10296
rect 1546 10240 1551 10296
rect 0 10238 1551 10240
rect 0 10208 800 10238
rect 1485 10235 1551 10238
rect 4317 9824 4637 9825
rect 4317 9760 4325 9824
rect 4389 9760 4405 9824
rect 4469 9760 4485 9824
rect 4549 9760 4565 9824
rect 4629 9760 4637 9824
rect 4317 9759 4637 9760
rect 7690 9824 8010 9825
rect 7690 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7938 9824
rect 8002 9760 8010 9824
rect 7690 9759 8010 9760
rect 2630 9280 2950 9281
rect 2630 9216 2638 9280
rect 2702 9216 2718 9280
rect 2782 9216 2798 9280
rect 2862 9216 2878 9280
rect 2942 9216 2950 9280
rect 2630 9215 2950 9216
rect 6004 9280 6324 9281
rect 6004 9216 6012 9280
rect 6076 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6324 9280
rect 6004 9215 6324 9216
rect 9377 9280 9697 9281
rect 9377 9216 9385 9280
rect 9449 9216 9465 9280
rect 9529 9216 9545 9280
rect 9609 9216 9625 9280
rect 9689 9216 9697 9280
rect 9377 9215 9697 9216
rect 4317 8736 4637 8737
rect 4317 8672 4325 8736
rect 4389 8672 4405 8736
rect 4469 8672 4485 8736
rect 4549 8672 4565 8736
rect 4629 8672 4637 8736
rect 4317 8671 4637 8672
rect 7690 8736 8010 8737
rect 7690 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7938 8736
rect 8002 8672 8010 8736
rect 7690 8671 8010 8672
rect 2630 8192 2950 8193
rect 2630 8128 2638 8192
rect 2702 8128 2718 8192
rect 2782 8128 2798 8192
rect 2862 8128 2878 8192
rect 2942 8128 2950 8192
rect 2630 8127 2950 8128
rect 6004 8192 6324 8193
rect 6004 8128 6012 8192
rect 6076 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6324 8192
rect 6004 8127 6324 8128
rect 9377 8192 9697 8193
rect 9377 8128 9385 8192
rect 9449 8128 9465 8192
rect 9529 8128 9545 8192
rect 9609 8128 9625 8192
rect 9689 8128 9697 8192
rect 9377 8127 9697 8128
rect 4317 7648 4637 7649
rect 4317 7584 4325 7648
rect 4389 7584 4405 7648
rect 4469 7584 4485 7648
rect 4549 7584 4565 7648
rect 4629 7584 4637 7648
rect 4317 7583 4637 7584
rect 7690 7648 8010 7649
rect 7690 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7938 7648
rect 8002 7584 8010 7648
rect 7690 7583 8010 7584
rect 10409 7578 10475 7581
rect 11529 7578 12329 7608
rect 10409 7576 12329 7578
rect 10409 7520 10414 7576
rect 10470 7520 12329 7576
rect 10409 7518 12329 7520
rect 10409 7515 10475 7518
rect 11529 7488 12329 7518
rect 2630 7104 2950 7105
rect 2630 7040 2638 7104
rect 2702 7040 2718 7104
rect 2782 7040 2798 7104
rect 2862 7040 2878 7104
rect 2942 7040 2950 7104
rect 2630 7039 2950 7040
rect 6004 7104 6324 7105
rect 6004 7040 6012 7104
rect 6076 7040 6092 7104
rect 6156 7040 6172 7104
rect 6236 7040 6252 7104
rect 6316 7040 6324 7104
rect 6004 7039 6324 7040
rect 9377 7104 9697 7105
rect 9377 7040 9385 7104
rect 9449 7040 9465 7104
rect 9529 7040 9545 7104
rect 9609 7040 9625 7104
rect 9689 7040 9697 7104
rect 9377 7039 9697 7040
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 4317 6560 4637 6561
rect 4317 6496 4325 6560
rect 4389 6496 4405 6560
rect 4469 6496 4485 6560
rect 4549 6496 4565 6560
rect 4629 6496 4637 6560
rect 4317 6495 4637 6496
rect 7690 6560 8010 6561
rect 7690 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7938 6560
rect 8002 6496 8010 6560
rect 7690 6495 8010 6496
rect 2630 6016 2950 6017
rect 2630 5952 2638 6016
rect 2702 5952 2718 6016
rect 2782 5952 2798 6016
rect 2862 5952 2878 6016
rect 2942 5952 2950 6016
rect 2630 5951 2950 5952
rect 6004 6016 6324 6017
rect 6004 5952 6012 6016
rect 6076 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6324 6016
rect 6004 5951 6324 5952
rect 9377 6016 9697 6017
rect 9377 5952 9385 6016
rect 9449 5952 9465 6016
rect 9529 5952 9545 6016
rect 9609 5952 9625 6016
rect 9689 5952 9697 6016
rect 9377 5951 9697 5952
rect 4317 5472 4637 5473
rect 4317 5408 4325 5472
rect 4389 5408 4405 5472
rect 4469 5408 4485 5472
rect 4549 5408 4565 5472
rect 4629 5408 4637 5472
rect 4317 5407 4637 5408
rect 7690 5472 8010 5473
rect 7690 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7938 5472
rect 8002 5408 8010 5472
rect 7690 5407 8010 5408
rect 2630 4928 2950 4929
rect 2630 4864 2638 4928
rect 2702 4864 2718 4928
rect 2782 4864 2798 4928
rect 2862 4864 2878 4928
rect 2942 4864 2950 4928
rect 2630 4863 2950 4864
rect 6004 4928 6324 4929
rect 6004 4864 6012 4928
rect 6076 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6324 4928
rect 6004 4863 6324 4864
rect 9377 4928 9697 4929
rect 9377 4864 9385 4928
rect 9449 4864 9465 4928
rect 9529 4864 9545 4928
rect 9609 4864 9625 4928
rect 9689 4864 9697 4928
rect 9377 4863 9697 4864
rect 4317 4384 4637 4385
rect 4317 4320 4325 4384
rect 4389 4320 4405 4384
rect 4469 4320 4485 4384
rect 4549 4320 4565 4384
rect 4629 4320 4637 4384
rect 4317 4319 4637 4320
rect 7690 4384 8010 4385
rect 7690 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7938 4384
rect 8002 4320 8010 4384
rect 7690 4319 8010 4320
rect 10501 4178 10567 4181
rect 11529 4178 12329 4208
rect 10501 4176 12329 4178
rect 10501 4120 10506 4176
rect 10562 4120 12329 4176
rect 10501 4118 12329 4120
rect 10501 4115 10567 4118
rect 11529 4088 12329 4118
rect 2630 3840 2950 3841
rect 2630 3776 2638 3840
rect 2702 3776 2718 3840
rect 2782 3776 2798 3840
rect 2862 3776 2878 3840
rect 2942 3776 2950 3840
rect 2630 3775 2950 3776
rect 6004 3840 6324 3841
rect 6004 3776 6012 3840
rect 6076 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6324 3840
rect 6004 3775 6324 3776
rect 9377 3840 9697 3841
rect 9377 3776 9385 3840
rect 9449 3776 9465 3840
rect 9529 3776 9545 3840
rect 9609 3776 9625 3840
rect 9689 3776 9697 3840
rect 9377 3775 9697 3776
rect 0 3498 800 3528
rect 1485 3498 1551 3501
rect 0 3496 1551 3498
rect 0 3440 1490 3496
rect 1546 3440 1551 3496
rect 0 3438 1551 3440
rect 0 3408 800 3438
rect 1485 3435 1551 3438
rect 4317 3296 4637 3297
rect 4317 3232 4325 3296
rect 4389 3232 4405 3296
rect 4469 3232 4485 3296
rect 4549 3232 4565 3296
rect 4629 3232 4637 3296
rect 4317 3231 4637 3232
rect 7690 3296 8010 3297
rect 7690 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7938 3296
rect 8002 3232 8010 3296
rect 7690 3231 8010 3232
rect 2630 2752 2950 2753
rect 2630 2688 2638 2752
rect 2702 2688 2718 2752
rect 2782 2688 2798 2752
rect 2862 2688 2878 2752
rect 2942 2688 2950 2752
rect 2630 2687 2950 2688
rect 6004 2752 6324 2753
rect 6004 2688 6012 2752
rect 6076 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6324 2752
rect 6004 2687 6324 2688
rect 9377 2752 9697 2753
rect 9377 2688 9385 2752
rect 9449 2688 9465 2752
rect 9529 2688 9545 2752
rect 9609 2688 9625 2752
rect 9689 2688 9697 2752
rect 9377 2687 9697 2688
rect 4317 2208 4637 2209
rect 4317 2144 4325 2208
rect 4389 2144 4405 2208
rect 4469 2144 4485 2208
rect 4549 2144 4565 2208
rect 4629 2144 4637 2208
rect 4317 2143 4637 2144
rect 7690 2208 8010 2209
rect 7690 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7938 2208
rect 8002 2144 8010 2208
rect 7690 2143 8010 2144
rect 10409 778 10475 781
rect 11529 778 12329 808
rect 10409 776 12329 778
rect 10409 720 10414 776
rect 10470 720 12329 776
rect 10409 718 12329 720
rect 10409 715 10475 718
rect 11529 688 12329 718
<< via3 >>
rect 4325 11996 4389 12000
rect 4325 11940 4329 11996
rect 4329 11940 4385 11996
rect 4385 11940 4389 11996
rect 4325 11936 4389 11940
rect 4405 11996 4469 12000
rect 4405 11940 4409 11996
rect 4409 11940 4465 11996
rect 4465 11940 4469 11996
rect 4405 11936 4469 11940
rect 4485 11996 4549 12000
rect 4485 11940 4489 11996
rect 4489 11940 4545 11996
rect 4545 11940 4549 11996
rect 4485 11936 4549 11940
rect 4565 11996 4629 12000
rect 4565 11940 4569 11996
rect 4569 11940 4625 11996
rect 4625 11940 4629 11996
rect 4565 11936 4629 11940
rect 7698 11996 7762 12000
rect 7698 11940 7702 11996
rect 7702 11940 7758 11996
rect 7758 11940 7762 11996
rect 7698 11936 7762 11940
rect 7778 11996 7842 12000
rect 7778 11940 7782 11996
rect 7782 11940 7838 11996
rect 7838 11940 7842 11996
rect 7778 11936 7842 11940
rect 7858 11996 7922 12000
rect 7858 11940 7862 11996
rect 7862 11940 7918 11996
rect 7918 11940 7922 11996
rect 7858 11936 7922 11940
rect 7938 11996 8002 12000
rect 7938 11940 7942 11996
rect 7942 11940 7998 11996
rect 7998 11940 8002 11996
rect 7938 11936 8002 11940
rect 2638 11452 2702 11456
rect 2638 11396 2642 11452
rect 2642 11396 2698 11452
rect 2698 11396 2702 11452
rect 2638 11392 2702 11396
rect 2718 11452 2782 11456
rect 2718 11396 2722 11452
rect 2722 11396 2778 11452
rect 2778 11396 2782 11452
rect 2718 11392 2782 11396
rect 2798 11452 2862 11456
rect 2798 11396 2802 11452
rect 2802 11396 2858 11452
rect 2858 11396 2862 11452
rect 2798 11392 2862 11396
rect 2878 11452 2942 11456
rect 2878 11396 2882 11452
rect 2882 11396 2938 11452
rect 2938 11396 2942 11452
rect 2878 11392 2942 11396
rect 6012 11452 6076 11456
rect 6012 11396 6016 11452
rect 6016 11396 6072 11452
rect 6072 11396 6076 11452
rect 6012 11392 6076 11396
rect 6092 11452 6156 11456
rect 6092 11396 6096 11452
rect 6096 11396 6152 11452
rect 6152 11396 6156 11452
rect 6092 11392 6156 11396
rect 6172 11452 6236 11456
rect 6172 11396 6176 11452
rect 6176 11396 6232 11452
rect 6232 11396 6236 11452
rect 6172 11392 6236 11396
rect 6252 11452 6316 11456
rect 6252 11396 6256 11452
rect 6256 11396 6312 11452
rect 6312 11396 6316 11452
rect 6252 11392 6316 11396
rect 9385 11452 9449 11456
rect 9385 11396 9389 11452
rect 9389 11396 9445 11452
rect 9445 11396 9449 11452
rect 9385 11392 9449 11396
rect 9465 11452 9529 11456
rect 9465 11396 9469 11452
rect 9469 11396 9525 11452
rect 9525 11396 9529 11452
rect 9465 11392 9529 11396
rect 9545 11452 9609 11456
rect 9545 11396 9549 11452
rect 9549 11396 9605 11452
rect 9605 11396 9609 11452
rect 9545 11392 9609 11396
rect 9625 11452 9689 11456
rect 9625 11396 9629 11452
rect 9629 11396 9685 11452
rect 9685 11396 9689 11452
rect 9625 11392 9689 11396
rect 4325 10908 4389 10912
rect 4325 10852 4329 10908
rect 4329 10852 4385 10908
rect 4385 10852 4389 10908
rect 4325 10848 4389 10852
rect 4405 10908 4469 10912
rect 4405 10852 4409 10908
rect 4409 10852 4465 10908
rect 4465 10852 4469 10908
rect 4405 10848 4469 10852
rect 4485 10908 4549 10912
rect 4485 10852 4489 10908
rect 4489 10852 4545 10908
rect 4545 10852 4549 10908
rect 4485 10848 4549 10852
rect 4565 10908 4629 10912
rect 4565 10852 4569 10908
rect 4569 10852 4625 10908
rect 4625 10852 4629 10908
rect 4565 10848 4629 10852
rect 7698 10908 7762 10912
rect 7698 10852 7702 10908
rect 7702 10852 7758 10908
rect 7758 10852 7762 10908
rect 7698 10848 7762 10852
rect 7778 10908 7842 10912
rect 7778 10852 7782 10908
rect 7782 10852 7838 10908
rect 7838 10852 7842 10908
rect 7778 10848 7842 10852
rect 7858 10908 7922 10912
rect 7858 10852 7862 10908
rect 7862 10852 7918 10908
rect 7918 10852 7922 10908
rect 7858 10848 7922 10852
rect 7938 10908 8002 10912
rect 7938 10852 7942 10908
rect 7942 10852 7998 10908
rect 7998 10852 8002 10908
rect 7938 10848 8002 10852
rect 2638 10364 2702 10368
rect 2638 10308 2642 10364
rect 2642 10308 2698 10364
rect 2698 10308 2702 10364
rect 2638 10304 2702 10308
rect 2718 10364 2782 10368
rect 2718 10308 2722 10364
rect 2722 10308 2778 10364
rect 2778 10308 2782 10364
rect 2718 10304 2782 10308
rect 2798 10364 2862 10368
rect 2798 10308 2802 10364
rect 2802 10308 2858 10364
rect 2858 10308 2862 10364
rect 2798 10304 2862 10308
rect 2878 10364 2942 10368
rect 2878 10308 2882 10364
rect 2882 10308 2938 10364
rect 2938 10308 2942 10364
rect 2878 10304 2942 10308
rect 6012 10364 6076 10368
rect 6012 10308 6016 10364
rect 6016 10308 6072 10364
rect 6072 10308 6076 10364
rect 6012 10304 6076 10308
rect 6092 10364 6156 10368
rect 6092 10308 6096 10364
rect 6096 10308 6152 10364
rect 6152 10308 6156 10364
rect 6092 10304 6156 10308
rect 6172 10364 6236 10368
rect 6172 10308 6176 10364
rect 6176 10308 6232 10364
rect 6232 10308 6236 10364
rect 6172 10304 6236 10308
rect 6252 10364 6316 10368
rect 6252 10308 6256 10364
rect 6256 10308 6312 10364
rect 6312 10308 6316 10364
rect 6252 10304 6316 10308
rect 9385 10364 9449 10368
rect 9385 10308 9389 10364
rect 9389 10308 9445 10364
rect 9445 10308 9449 10364
rect 9385 10304 9449 10308
rect 9465 10364 9529 10368
rect 9465 10308 9469 10364
rect 9469 10308 9525 10364
rect 9525 10308 9529 10364
rect 9465 10304 9529 10308
rect 9545 10364 9609 10368
rect 9545 10308 9549 10364
rect 9549 10308 9605 10364
rect 9605 10308 9609 10364
rect 9545 10304 9609 10308
rect 9625 10364 9689 10368
rect 9625 10308 9629 10364
rect 9629 10308 9685 10364
rect 9685 10308 9689 10364
rect 9625 10304 9689 10308
rect 4325 9820 4389 9824
rect 4325 9764 4329 9820
rect 4329 9764 4385 9820
rect 4385 9764 4389 9820
rect 4325 9760 4389 9764
rect 4405 9820 4469 9824
rect 4405 9764 4409 9820
rect 4409 9764 4465 9820
rect 4465 9764 4469 9820
rect 4405 9760 4469 9764
rect 4485 9820 4549 9824
rect 4485 9764 4489 9820
rect 4489 9764 4545 9820
rect 4545 9764 4549 9820
rect 4485 9760 4549 9764
rect 4565 9820 4629 9824
rect 4565 9764 4569 9820
rect 4569 9764 4625 9820
rect 4625 9764 4629 9820
rect 4565 9760 4629 9764
rect 7698 9820 7762 9824
rect 7698 9764 7702 9820
rect 7702 9764 7758 9820
rect 7758 9764 7762 9820
rect 7698 9760 7762 9764
rect 7778 9820 7842 9824
rect 7778 9764 7782 9820
rect 7782 9764 7838 9820
rect 7838 9764 7842 9820
rect 7778 9760 7842 9764
rect 7858 9820 7922 9824
rect 7858 9764 7862 9820
rect 7862 9764 7918 9820
rect 7918 9764 7922 9820
rect 7858 9760 7922 9764
rect 7938 9820 8002 9824
rect 7938 9764 7942 9820
rect 7942 9764 7998 9820
rect 7998 9764 8002 9820
rect 7938 9760 8002 9764
rect 2638 9276 2702 9280
rect 2638 9220 2642 9276
rect 2642 9220 2698 9276
rect 2698 9220 2702 9276
rect 2638 9216 2702 9220
rect 2718 9276 2782 9280
rect 2718 9220 2722 9276
rect 2722 9220 2778 9276
rect 2778 9220 2782 9276
rect 2718 9216 2782 9220
rect 2798 9276 2862 9280
rect 2798 9220 2802 9276
rect 2802 9220 2858 9276
rect 2858 9220 2862 9276
rect 2798 9216 2862 9220
rect 2878 9276 2942 9280
rect 2878 9220 2882 9276
rect 2882 9220 2938 9276
rect 2938 9220 2942 9276
rect 2878 9216 2942 9220
rect 6012 9276 6076 9280
rect 6012 9220 6016 9276
rect 6016 9220 6072 9276
rect 6072 9220 6076 9276
rect 6012 9216 6076 9220
rect 6092 9276 6156 9280
rect 6092 9220 6096 9276
rect 6096 9220 6152 9276
rect 6152 9220 6156 9276
rect 6092 9216 6156 9220
rect 6172 9276 6236 9280
rect 6172 9220 6176 9276
rect 6176 9220 6232 9276
rect 6232 9220 6236 9276
rect 6172 9216 6236 9220
rect 6252 9276 6316 9280
rect 6252 9220 6256 9276
rect 6256 9220 6312 9276
rect 6312 9220 6316 9276
rect 6252 9216 6316 9220
rect 9385 9276 9449 9280
rect 9385 9220 9389 9276
rect 9389 9220 9445 9276
rect 9445 9220 9449 9276
rect 9385 9216 9449 9220
rect 9465 9276 9529 9280
rect 9465 9220 9469 9276
rect 9469 9220 9525 9276
rect 9525 9220 9529 9276
rect 9465 9216 9529 9220
rect 9545 9276 9609 9280
rect 9545 9220 9549 9276
rect 9549 9220 9605 9276
rect 9605 9220 9609 9276
rect 9545 9216 9609 9220
rect 9625 9276 9689 9280
rect 9625 9220 9629 9276
rect 9629 9220 9685 9276
rect 9685 9220 9689 9276
rect 9625 9216 9689 9220
rect 4325 8732 4389 8736
rect 4325 8676 4329 8732
rect 4329 8676 4385 8732
rect 4385 8676 4389 8732
rect 4325 8672 4389 8676
rect 4405 8732 4469 8736
rect 4405 8676 4409 8732
rect 4409 8676 4465 8732
rect 4465 8676 4469 8732
rect 4405 8672 4469 8676
rect 4485 8732 4549 8736
rect 4485 8676 4489 8732
rect 4489 8676 4545 8732
rect 4545 8676 4549 8732
rect 4485 8672 4549 8676
rect 4565 8732 4629 8736
rect 4565 8676 4569 8732
rect 4569 8676 4625 8732
rect 4625 8676 4629 8732
rect 4565 8672 4629 8676
rect 7698 8732 7762 8736
rect 7698 8676 7702 8732
rect 7702 8676 7758 8732
rect 7758 8676 7762 8732
rect 7698 8672 7762 8676
rect 7778 8732 7842 8736
rect 7778 8676 7782 8732
rect 7782 8676 7838 8732
rect 7838 8676 7842 8732
rect 7778 8672 7842 8676
rect 7858 8732 7922 8736
rect 7858 8676 7862 8732
rect 7862 8676 7918 8732
rect 7918 8676 7922 8732
rect 7858 8672 7922 8676
rect 7938 8732 8002 8736
rect 7938 8676 7942 8732
rect 7942 8676 7998 8732
rect 7998 8676 8002 8732
rect 7938 8672 8002 8676
rect 2638 8188 2702 8192
rect 2638 8132 2642 8188
rect 2642 8132 2698 8188
rect 2698 8132 2702 8188
rect 2638 8128 2702 8132
rect 2718 8188 2782 8192
rect 2718 8132 2722 8188
rect 2722 8132 2778 8188
rect 2778 8132 2782 8188
rect 2718 8128 2782 8132
rect 2798 8188 2862 8192
rect 2798 8132 2802 8188
rect 2802 8132 2858 8188
rect 2858 8132 2862 8188
rect 2798 8128 2862 8132
rect 2878 8188 2942 8192
rect 2878 8132 2882 8188
rect 2882 8132 2938 8188
rect 2938 8132 2942 8188
rect 2878 8128 2942 8132
rect 6012 8188 6076 8192
rect 6012 8132 6016 8188
rect 6016 8132 6072 8188
rect 6072 8132 6076 8188
rect 6012 8128 6076 8132
rect 6092 8188 6156 8192
rect 6092 8132 6096 8188
rect 6096 8132 6152 8188
rect 6152 8132 6156 8188
rect 6092 8128 6156 8132
rect 6172 8188 6236 8192
rect 6172 8132 6176 8188
rect 6176 8132 6232 8188
rect 6232 8132 6236 8188
rect 6172 8128 6236 8132
rect 6252 8188 6316 8192
rect 6252 8132 6256 8188
rect 6256 8132 6312 8188
rect 6312 8132 6316 8188
rect 6252 8128 6316 8132
rect 9385 8188 9449 8192
rect 9385 8132 9389 8188
rect 9389 8132 9445 8188
rect 9445 8132 9449 8188
rect 9385 8128 9449 8132
rect 9465 8188 9529 8192
rect 9465 8132 9469 8188
rect 9469 8132 9525 8188
rect 9525 8132 9529 8188
rect 9465 8128 9529 8132
rect 9545 8188 9609 8192
rect 9545 8132 9549 8188
rect 9549 8132 9605 8188
rect 9605 8132 9609 8188
rect 9545 8128 9609 8132
rect 9625 8188 9689 8192
rect 9625 8132 9629 8188
rect 9629 8132 9685 8188
rect 9685 8132 9689 8188
rect 9625 8128 9689 8132
rect 4325 7644 4389 7648
rect 4325 7588 4329 7644
rect 4329 7588 4385 7644
rect 4385 7588 4389 7644
rect 4325 7584 4389 7588
rect 4405 7644 4469 7648
rect 4405 7588 4409 7644
rect 4409 7588 4465 7644
rect 4465 7588 4469 7644
rect 4405 7584 4469 7588
rect 4485 7644 4549 7648
rect 4485 7588 4489 7644
rect 4489 7588 4545 7644
rect 4545 7588 4549 7644
rect 4485 7584 4549 7588
rect 4565 7644 4629 7648
rect 4565 7588 4569 7644
rect 4569 7588 4625 7644
rect 4625 7588 4629 7644
rect 4565 7584 4629 7588
rect 7698 7644 7762 7648
rect 7698 7588 7702 7644
rect 7702 7588 7758 7644
rect 7758 7588 7762 7644
rect 7698 7584 7762 7588
rect 7778 7644 7842 7648
rect 7778 7588 7782 7644
rect 7782 7588 7838 7644
rect 7838 7588 7842 7644
rect 7778 7584 7842 7588
rect 7858 7644 7922 7648
rect 7858 7588 7862 7644
rect 7862 7588 7918 7644
rect 7918 7588 7922 7644
rect 7858 7584 7922 7588
rect 7938 7644 8002 7648
rect 7938 7588 7942 7644
rect 7942 7588 7998 7644
rect 7998 7588 8002 7644
rect 7938 7584 8002 7588
rect 2638 7100 2702 7104
rect 2638 7044 2642 7100
rect 2642 7044 2698 7100
rect 2698 7044 2702 7100
rect 2638 7040 2702 7044
rect 2718 7100 2782 7104
rect 2718 7044 2722 7100
rect 2722 7044 2778 7100
rect 2778 7044 2782 7100
rect 2718 7040 2782 7044
rect 2798 7100 2862 7104
rect 2798 7044 2802 7100
rect 2802 7044 2858 7100
rect 2858 7044 2862 7100
rect 2798 7040 2862 7044
rect 2878 7100 2942 7104
rect 2878 7044 2882 7100
rect 2882 7044 2938 7100
rect 2938 7044 2942 7100
rect 2878 7040 2942 7044
rect 6012 7100 6076 7104
rect 6012 7044 6016 7100
rect 6016 7044 6072 7100
rect 6072 7044 6076 7100
rect 6012 7040 6076 7044
rect 6092 7100 6156 7104
rect 6092 7044 6096 7100
rect 6096 7044 6152 7100
rect 6152 7044 6156 7100
rect 6092 7040 6156 7044
rect 6172 7100 6236 7104
rect 6172 7044 6176 7100
rect 6176 7044 6232 7100
rect 6232 7044 6236 7100
rect 6172 7040 6236 7044
rect 6252 7100 6316 7104
rect 6252 7044 6256 7100
rect 6256 7044 6312 7100
rect 6312 7044 6316 7100
rect 6252 7040 6316 7044
rect 9385 7100 9449 7104
rect 9385 7044 9389 7100
rect 9389 7044 9445 7100
rect 9445 7044 9449 7100
rect 9385 7040 9449 7044
rect 9465 7100 9529 7104
rect 9465 7044 9469 7100
rect 9469 7044 9525 7100
rect 9525 7044 9529 7100
rect 9465 7040 9529 7044
rect 9545 7100 9609 7104
rect 9545 7044 9549 7100
rect 9549 7044 9605 7100
rect 9605 7044 9609 7100
rect 9545 7040 9609 7044
rect 9625 7100 9689 7104
rect 9625 7044 9629 7100
rect 9629 7044 9685 7100
rect 9685 7044 9689 7100
rect 9625 7040 9689 7044
rect 4325 6556 4389 6560
rect 4325 6500 4329 6556
rect 4329 6500 4385 6556
rect 4385 6500 4389 6556
rect 4325 6496 4389 6500
rect 4405 6556 4469 6560
rect 4405 6500 4409 6556
rect 4409 6500 4465 6556
rect 4465 6500 4469 6556
rect 4405 6496 4469 6500
rect 4485 6556 4549 6560
rect 4485 6500 4489 6556
rect 4489 6500 4545 6556
rect 4545 6500 4549 6556
rect 4485 6496 4549 6500
rect 4565 6556 4629 6560
rect 4565 6500 4569 6556
rect 4569 6500 4625 6556
rect 4625 6500 4629 6556
rect 4565 6496 4629 6500
rect 7698 6556 7762 6560
rect 7698 6500 7702 6556
rect 7702 6500 7758 6556
rect 7758 6500 7762 6556
rect 7698 6496 7762 6500
rect 7778 6556 7842 6560
rect 7778 6500 7782 6556
rect 7782 6500 7838 6556
rect 7838 6500 7842 6556
rect 7778 6496 7842 6500
rect 7858 6556 7922 6560
rect 7858 6500 7862 6556
rect 7862 6500 7918 6556
rect 7918 6500 7922 6556
rect 7858 6496 7922 6500
rect 7938 6556 8002 6560
rect 7938 6500 7942 6556
rect 7942 6500 7998 6556
rect 7998 6500 8002 6556
rect 7938 6496 8002 6500
rect 2638 6012 2702 6016
rect 2638 5956 2642 6012
rect 2642 5956 2698 6012
rect 2698 5956 2702 6012
rect 2638 5952 2702 5956
rect 2718 6012 2782 6016
rect 2718 5956 2722 6012
rect 2722 5956 2778 6012
rect 2778 5956 2782 6012
rect 2718 5952 2782 5956
rect 2798 6012 2862 6016
rect 2798 5956 2802 6012
rect 2802 5956 2858 6012
rect 2858 5956 2862 6012
rect 2798 5952 2862 5956
rect 2878 6012 2942 6016
rect 2878 5956 2882 6012
rect 2882 5956 2938 6012
rect 2938 5956 2942 6012
rect 2878 5952 2942 5956
rect 6012 6012 6076 6016
rect 6012 5956 6016 6012
rect 6016 5956 6072 6012
rect 6072 5956 6076 6012
rect 6012 5952 6076 5956
rect 6092 6012 6156 6016
rect 6092 5956 6096 6012
rect 6096 5956 6152 6012
rect 6152 5956 6156 6012
rect 6092 5952 6156 5956
rect 6172 6012 6236 6016
rect 6172 5956 6176 6012
rect 6176 5956 6232 6012
rect 6232 5956 6236 6012
rect 6172 5952 6236 5956
rect 6252 6012 6316 6016
rect 6252 5956 6256 6012
rect 6256 5956 6312 6012
rect 6312 5956 6316 6012
rect 6252 5952 6316 5956
rect 9385 6012 9449 6016
rect 9385 5956 9389 6012
rect 9389 5956 9445 6012
rect 9445 5956 9449 6012
rect 9385 5952 9449 5956
rect 9465 6012 9529 6016
rect 9465 5956 9469 6012
rect 9469 5956 9525 6012
rect 9525 5956 9529 6012
rect 9465 5952 9529 5956
rect 9545 6012 9609 6016
rect 9545 5956 9549 6012
rect 9549 5956 9605 6012
rect 9605 5956 9609 6012
rect 9545 5952 9609 5956
rect 9625 6012 9689 6016
rect 9625 5956 9629 6012
rect 9629 5956 9685 6012
rect 9685 5956 9689 6012
rect 9625 5952 9689 5956
rect 4325 5468 4389 5472
rect 4325 5412 4329 5468
rect 4329 5412 4385 5468
rect 4385 5412 4389 5468
rect 4325 5408 4389 5412
rect 4405 5468 4469 5472
rect 4405 5412 4409 5468
rect 4409 5412 4465 5468
rect 4465 5412 4469 5468
rect 4405 5408 4469 5412
rect 4485 5468 4549 5472
rect 4485 5412 4489 5468
rect 4489 5412 4545 5468
rect 4545 5412 4549 5468
rect 4485 5408 4549 5412
rect 4565 5468 4629 5472
rect 4565 5412 4569 5468
rect 4569 5412 4625 5468
rect 4625 5412 4629 5468
rect 4565 5408 4629 5412
rect 7698 5468 7762 5472
rect 7698 5412 7702 5468
rect 7702 5412 7758 5468
rect 7758 5412 7762 5468
rect 7698 5408 7762 5412
rect 7778 5468 7842 5472
rect 7778 5412 7782 5468
rect 7782 5412 7838 5468
rect 7838 5412 7842 5468
rect 7778 5408 7842 5412
rect 7858 5468 7922 5472
rect 7858 5412 7862 5468
rect 7862 5412 7918 5468
rect 7918 5412 7922 5468
rect 7858 5408 7922 5412
rect 7938 5468 8002 5472
rect 7938 5412 7942 5468
rect 7942 5412 7998 5468
rect 7998 5412 8002 5468
rect 7938 5408 8002 5412
rect 2638 4924 2702 4928
rect 2638 4868 2642 4924
rect 2642 4868 2698 4924
rect 2698 4868 2702 4924
rect 2638 4864 2702 4868
rect 2718 4924 2782 4928
rect 2718 4868 2722 4924
rect 2722 4868 2778 4924
rect 2778 4868 2782 4924
rect 2718 4864 2782 4868
rect 2798 4924 2862 4928
rect 2798 4868 2802 4924
rect 2802 4868 2858 4924
rect 2858 4868 2862 4924
rect 2798 4864 2862 4868
rect 2878 4924 2942 4928
rect 2878 4868 2882 4924
rect 2882 4868 2938 4924
rect 2938 4868 2942 4924
rect 2878 4864 2942 4868
rect 6012 4924 6076 4928
rect 6012 4868 6016 4924
rect 6016 4868 6072 4924
rect 6072 4868 6076 4924
rect 6012 4864 6076 4868
rect 6092 4924 6156 4928
rect 6092 4868 6096 4924
rect 6096 4868 6152 4924
rect 6152 4868 6156 4924
rect 6092 4864 6156 4868
rect 6172 4924 6236 4928
rect 6172 4868 6176 4924
rect 6176 4868 6232 4924
rect 6232 4868 6236 4924
rect 6172 4864 6236 4868
rect 6252 4924 6316 4928
rect 6252 4868 6256 4924
rect 6256 4868 6312 4924
rect 6312 4868 6316 4924
rect 6252 4864 6316 4868
rect 9385 4924 9449 4928
rect 9385 4868 9389 4924
rect 9389 4868 9445 4924
rect 9445 4868 9449 4924
rect 9385 4864 9449 4868
rect 9465 4924 9529 4928
rect 9465 4868 9469 4924
rect 9469 4868 9525 4924
rect 9525 4868 9529 4924
rect 9465 4864 9529 4868
rect 9545 4924 9609 4928
rect 9545 4868 9549 4924
rect 9549 4868 9605 4924
rect 9605 4868 9609 4924
rect 9545 4864 9609 4868
rect 9625 4924 9689 4928
rect 9625 4868 9629 4924
rect 9629 4868 9685 4924
rect 9685 4868 9689 4924
rect 9625 4864 9689 4868
rect 4325 4380 4389 4384
rect 4325 4324 4329 4380
rect 4329 4324 4385 4380
rect 4385 4324 4389 4380
rect 4325 4320 4389 4324
rect 4405 4380 4469 4384
rect 4405 4324 4409 4380
rect 4409 4324 4465 4380
rect 4465 4324 4469 4380
rect 4405 4320 4469 4324
rect 4485 4380 4549 4384
rect 4485 4324 4489 4380
rect 4489 4324 4545 4380
rect 4545 4324 4549 4380
rect 4485 4320 4549 4324
rect 4565 4380 4629 4384
rect 4565 4324 4569 4380
rect 4569 4324 4625 4380
rect 4625 4324 4629 4380
rect 4565 4320 4629 4324
rect 7698 4380 7762 4384
rect 7698 4324 7702 4380
rect 7702 4324 7758 4380
rect 7758 4324 7762 4380
rect 7698 4320 7762 4324
rect 7778 4380 7842 4384
rect 7778 4324 7782 4380
rect 7782 4324 7838 4380
rect 7838 4324 7842 4380
rect 7778 4320 7842 4324
rect 7858 4380 7922 4384
rect 7858 4324 7862 4380
rect 7862 4324 7918 4380
rect 7918 4324 7922 4380
rect 7858 4320 7922 4324
rect 7938 4380 8002 4384
rect 7938 4324 7942 4380
rect 7942 4324 7998 4380
rect 7998 4324 8002 4380
rect 7938 4320 8002 4324
rect 2638 3836 2702 3840
rect 2638 3780 2642 3836
rect 2642 3780 2698 3836
rect 2698 3780 2702 3836
rect 2638 3776 2702 3780
rect 2718 3836 2782 3840
rect 2718 3780 2722 3836
rect 2722 3780 2778 3836
rect 2778 3780 2782 3836
rect 2718 3776 2782 3780
rect 2798 3836 2862 3840
rect 2798 3780 2802 3836
rect 2802 3780 2858 3836
rect 2858 3780 2862 3836
rect 2798 3776 2862 3780
rect 2878 3836 2942 3840
rect 2878 3780 2882 3836
rect 2882 3780 2938 3836
rect 2938 3780 2942 3836
rect 2878 3776 2942 3780
rect 6012 3836 6076 3840
rect 6012 3780 6016 3836
rect 6016 3780 6072 3836
rect 6072 3780 6076 3836
rect 6012 3776 6076 3780
rect 6092 3836 6156 3840
rect 6092 3780 6096 3836
rect 6096 3780 6152 3836
rect 6152 3780 6156 3836
rect 6092 3776 6156 3780
rect 6172 3836 6236 3840
rect 6172 3780 6176 3836
rect 6176 3780 6232 3836
rect 6232 3780 6236 3836
rect 6172 3776 6236 3780
rect 6252 3836 6316 3840
rect 6252 3780 6256 3836
rect 6256 3780 6312 3836
rect 6312 3780 6316 3836
rect 6252 3776 6316 3780
rect 9385 3836 9449 3840
rect 9385 3780 9389 3836
rect 9389 3780 9445 3836
rect 9445 3780 9449 3836
rect 9385 3776 9449 3780
rect 9465 3836 9529 3840
rect 9465 3780 9469 3836
rect 9469 3780 9525 3836
rect 9525 3780 9529 3836
rect 9465 3776 9529 3780
rect 9545 3836 9609 3840
rect 9545 3780 9549 3836
rect 9549 3780 9605 3836
rect 9605 3780 9609 3836
rect 9545 3776 9609 3780
rect 9625 3836 9689 3840
rect 9625 3780 9629 3836
rect 9629 3780 9685 3836
rect 9685 3780 9689 3836
rect 9625 3776 9689 3780
rect 4325 3292 4389 3296
rect 4325 3236 4329 3292
rect 4329 3236 4385 3292
rect 4385 3236 4389 3292
rect 4325 3232 4389 3236
rect 4405 3292 4469 3296
rect 4405 3236 4409 3292
rect 4409 3236 4465 3292
rect 4465 3236 4469 3292
rect 4405 3232 4469 3236
rect 4485 3292 4549 3296
rect 4485 3236 4489 3292
rect 4489 3236 4545 3292
rect 4545 3236 4549 3292
rect 4485 3232 4549 3236
rect 4565 3292 4629 3296
rect 4565 3236 4569 3292
rect 4569 3236 4625 3292
rect 4625 3236 4629 3292
rect 4565 3232 4629 3236
rect 7698 3292 7762 3296
rect 7698 3236 7702 3292
rect 7702 3236 7758 3292
rect 7758 3236 7762 3292
rect 7698 3232 7762 3236
rect 7778 3292 7842 3296
rect 7778 3236 7782 3292
rect 7782 3236 7838 3292
rect 7838 3236 7842 3292
rect 7778 3232 7842 3236
rect 7858 3292 7922 3296
rect 7858 3236 7862 3292
rect 7862 3236 7918 3292
rect 7918 3236 7922 3292
rect 7858 3232 7922 3236
rect 7938 3292 8002 3296
rect 7938 3236 7942 3292
rect 7942 3236 7998 3292
rect 7998 3236 8002 3292
rect 7938 3232 8002 3236
rect 2638 2748 2702 2752
rect 2638 2692 2642 2748
rect 2642 2692 2698 2748
rect 2698 2692 2702 2748
rect 2638 2688 2702 2692
rect 2718 2748 2782 2752
rect 2718 2692 2722 2748
rect 2722 2692 2778 2748
rect 2778 2692 2782 2748
rect 2718 2688 2782 2692
rect 2798 2748 2862 2752
rect 2798 2692 2802 2748
rect 2802 2692 2858 2748
rect 2858 2692 2862 2748
rect 2798 2688 2862 2692
rect 2878 2748 2942 2752
rect 2878 2692 2882 2748
rect 2882 2692 2938 2748
rect 2938 2692 2942 2748
rect 2878 2688 2942 2692
rect 6012 2748 6076 2752
rect 6012 2692 6016 2748
rect 6016 2692 6072 2748
rect 6072 2692 6076 2748
rect 6012 2688 6076 2692
rect 6092 2748 6156 2752
rect 6092 2692 6096 2748
rect 6096 2692 6152 2748
rect 6152 2692 6156 2748
rect 6092 2688 6156 2692
rect 6172 2748 6236 2752
rect 6172 2692 6176 2748
rect 6176 2692 6232 2748
rect 6232 2692 6236 2748
rect 6172 2688 6236 2692
rect 6252 2748 6316 2752
rect 6252 2692 6256 2748
rect 6256 2692 6312 2748
rect 6312 2692 6316 2748
rect 6252 2688 6316 2692
rect 9385 2748 9449 2752
rect 9385 2692 9389 2748
rect 9389 2692 9445 2748
rect 9445 2692 9449 2748
rect 9385 2688 9449 2692
rect 9465 2748 9529 2752
rect 9465 2692 9469 2748
rect 9469 2692 9525 2748
rect 9525 2692 9529 2748
rect 9465 2688 9529 2692
rect 9545 2748 9609 2752
rect 9545 2692 9549 2748
rect 9549 2692 9605 2748
rect 9605 2692 9609 2748
rect 9545 2688 9609 2692
rect 9625 2748 9689 2752
rect 9625 2692 9629 2748
rect 9629 2692 9685 2748
rect 9685 2692 9689 2748
rect 9625 2688 9689 2692
rect 4325 2204 4389 2208
rect 4325 2148 4329 2204
rect 4329 2148 4385 2204
rect 4385 2148 4389 2204
rect 4325 2144 4389 2148
rect 4405 2204 4469 2208
rect 4405 2148 4409 2204
rect 4409 2148 4465 2204
rect 4465 2148 4469 2204
rect 4405 2144 4469 2148
rect 4485 2204 4549 2208
rect 4485 2148 4489 2204
rect 4489 2148 4545 2204
rect 4545 2148 4549 2204
rect 4485 2144 4549 2148
rect 4565 2204 4629 2208
rect 4565 2148 4569 2204
rect 4569 2148 4625 2204
rect 4625 2148 4629 2204
rect 4565 2144 4629 2148
rect 7698 2204 7762 2208
rect 7698 2148 7702 2204
rect 7702 2148 7758 2204
rect 7758 2148 7762 2204
rect 7698 2144 7762 2148
rect 7778 2204 7842 2208
rect 7778 2148 7782 2204
rect 7782 2148 7838 2204
rect 7838 2148 7842 2204
rect 7778 2144 7842 2148
rect 7858 2204 7922 2208
rect 7858 2148 7862 2204
rect 7862 2148 7918 2204
rect 7918 2148 7922 2204
rect 7858 2144 7922 2148
rect 7938 2204 8002 2208
rect 7938 2148 7942 2204
rect 7942 2148 7998 2204
rect 7998 2148 8002 2204
rect 7938 2144 8002 2148
<< metal4 >>
rect 2630 11456 2950 12016
rect 2630 11392 2638 11456
rect 2702 11392 2718 11456
rect 2782 11392 2798 11456
rect 2862 11392 2878 11456
rect 2942 11392 2950 11456
rect 2630 10406 2950 11392
rect 2630 10368 2672 10406
rect 2908 10368 2950 10406
rect 2630 10304 2638 10368
rect 2942 10304 2950 10368
rect 2630 10170 2672 10304
rect 2908 10170 2950 10304
rect 2630 9280 2950 10170
rect 2630 9216 2638 9280
rect 2702 9216 2718 9280
rect 2782 9216 2798 9280
rect 2862 9216 2878 9280
rect 2942 9216 2950 9280
rect 2630 8192 2950 9216
rect 2630 8128 2638 8192
rect 2702 8128 2718 8192
rect 2782 8128 2798 8192
rect 2862 8128 2878 8192
rect 2942 8128 2950 8192
rect 2630 7142 2950 8128
rect 2630 7104 2672 7142
rect 2908 7104 2950 7142
rect 2630 7040 2638 7104
rect 2942 7040 2950 7104
rect 2630 6906 2672 7040
rect 2908 6906 2950 7040
rect 2630 6016 2950 6906
rect 2630 5952 2638 6016
rect 2702 5952 2718 6016
rect 2782 5952 2798 6016
rect 2862 5952 2878 6016
rect 2942 5952 2950 6016
rect 2630 4928 2950 5952
rect 2630 4864 2638 4928
rect 2702 4864 2718 4928
rect 2782 4864 2798 4928
rect 2862 4864 2878 4928
rect 2942 4864 2950 4928
rect 2630 3878 2950 4864
rect 2630 3840 2672 3878
rect 2908 3840 2950 3878
rect 2630 3776 2638 3840
rect 2942 3776 2950 3840
rect 2630 3642 2672 3776
rect 2908 3642 2950 3776
rect 2630 2752 2950 3642
rect 2630 2688 2638 2752
rect 2702 2688 2718 2752
rect 2782 2688 2798 2752
rect 2862 2688 2878 2752
rect 2942 2688 2950 2752
rect 2630 2128 2950 2688
rect 4317 12000 4638 12016
rect 4317 11936 4325 12000
rect 4389 11936 4405 12000
rect 4469 11936 4485 12000
rect 4549 11936 4565 12000
rect 4629 11936 4638 12000
rect 4317 10912 4638 11936
rect 4317 10848 4325 10912
rect 4389 10848 4405 10912
rect 4469 10848 4485 10912
rect 4549 10848 4565 10912
rect 4629 10848 4638 10912
rect 4317 9824 4638 10848
rect 4317 9760 4325 9824
rect 4389 9760 4405 9824
rect 4469 9760 4485 9824
rect 4549 9760 4565 9824
rect 4629 9760 4638 9824
rect 4317 8774 4638 9760
rect 4317 8736 4359 8774
rect 4595 8736 4638 8774
rect 4317 8672 4325 8736
rect 4629 8672 4638 8736
rect 4317 8538 4359 8672
rect 4595 8538 4638 8672
rect 4317 7648 4638 8538
rect 4317 7584 4325 7648
rect 4389 7584 4405 7648
rect 4469 7584 4485 7648
rect 4549 7584 4565 7648
rect 4629 7584 4638 7648
rect 4317 6560 4638 7584
rect 4317 6496 4325 6560
rect 4389 6496 4405 6560
rect 4469 6496 4485 6560
rect 4549 6496 4565 6560
rect 4629 6496 4638 6560
rect 4317 5510 4638 6496
rect 4317 5472 4359 5510
rect 4595 5472 4638 5510
rect 4317 5408 4325 5472
rect 4629 5408 4638 5472
rect 4317 5274 4359 5408
rect 4595 5274 4638 5408
rect 4317 4384 4638 5274
rect 4317 4320 4325 4384
rect 4389 4320 4405 4384
rect 4469 4320 4485 4384
rect 4549 4320 4565 4384
rect 4629 4320 4638 4384
rect 4317 3296 4638 4320
rect 4317 3232 4325 3296
rect 4389 3232 4405 3296
rect 4469 3232 4485 3296
rect 4549 3232 4565 3296
rect 4629 3232 4638 3296
rect 4317 2208 4638 3232
rect 4317 2144 4325 2208
rect 4389 2144 4405 2208
rect 4469 2144 4485 2208
rect 4549 2144 4565 2208
rect 4629 2144 4638 2208
rect 4317 2128 4638 2144
rect 6004 11456 6324 12016
rect 6004 11392 6012 11456
rect 6076 11392 6092 11456
rect 6156 11392 6172 11456
rect 6236 11392 6252 11456
rect 6316 11392 6324 11456
rect 6004 10406 6324 11392
rect 6004 10368 6046 10406
rect 6282 10368 6324 10406
rect 6004 10304 6012 10368
rect 6316 10304 6324 10368
rect 6004 10170 6046 10304
rect 6282 10170 6324 10304
rect 6004 9280 6324 10170
rect 6004 9216 6012 9280
rect 6076 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6324 9280
rect 6004 8192 6324 9216
rect 6004 8128 6012 8192
rect 6076 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6324 8192
rect 6004 7142 6324 8128
rect 6004 7104 6046 7142
rect 6282 7104 6324 7142
rect 6004 7040 6012 7104
rect 6316 7040 6324 7104
rect 6004 6906 6046 7040
rect 6282 6906 6324 7040
rect 6004 6016 6324 6906
rect 6004 5952 6012 6016
rect 6076 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6324 6016
rect 6004 4928 6324 5952
rect 6004 4864 6012 4928
rect 6076 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6324 4928
rect 6004 3878 6324 4864
rect 6004 3840 6046 3878
rect 6282 3840 6324 3878
rect 6004 3776 6012 3840
rect 6316 3776 6324 3840
rect 6004 3642 6046 3776
rect 6282 3642 6324 3776
rect 6004 2752 6324 3642
rect 6004 2688 6012 2752
rect 6076 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6324 2752
rect 6004 2128 6324 2688
rect 7690 12000 8011 12016
rect 7690 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7938 12000
rect 8002 11936 8011 12000
rect 7690 10912 8011 11936
rect 7690 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7938 10912
rect 8002 10848 8011 10912
rect 7690 9824 8011 10848
rect 7690 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7938 9824
rect 8002 9760 8011 9824
rect 7690 8774 8011 9760
rect 7690 8736 7732 8774
rect 7968 8736 8011 8774
rect 7690 8672 7698 8736
rect 8002 8672 8011 8736
rect 7690 8538 7732 8672
rect 7968 8538 8011 8672
rect 7690 7648 8011 8538
rect 7690 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7938 7648
rect 8002 7584 8011 7648
rect 7690 6560 8011 7584
rect 7690 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7938 6560
rect 8002 6496 8011 6560
rect 7690 5510 8011 6496
rect 7690 5472 7732 5510
rect 7968 5472 8011 5510
rect 7690 5408 7698 5472
rect 8002 5408 8011 5472
rect 7690 5274 7732 5408
rect 7968 5274 8011 5408
rect 7690 4384 8011 5274
rect 7690 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7938 4384
rect 8002 4320 8011 4384
rect 7690 3296 8011 4320
rect 7690 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7938 3296
rect 8002 3232 8011 3296
rect 7690 2208 8011 3232
rect 7690 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7938 2208
rect 8002 2144 8011 2208
rect 7690 2128 8011 2144
rect 9377 11456 9697 12016
rect 9377 11392 9385 11456
rect 9449 11392 9465 11456
rect 9529 11392 9545 11456
rect 9609 11392 9625 11456
rect 9689 11392 9697 11456
rect 9377 10406 9697 11392
rect 9377 10368 9419 10406
rect 9655 10368 9697 10406
rect 9377 10304 9385 10368
rect 9689 10304 9697 10368
rect 9377 10170 9419 10304
rect 9655 10170 9697 10304
rect 9377 9280 9697 10170
rect 9377 9216 9385 9280
rect 9449 9216 9465 9280
rect 9529 9216 9545 9280
rect 9609 9216 9625 9280
rect 9689 9216 9697 9280
rect 9377 8192 9697 9216
rect 9377 8128 9385 8192
rect 9449 8128 9465 8192
rect 9529 8128 9545 8192
rect 9609 8128 9625 8192
rect 9689 8128 9697 8192
rect 9377 7142 9697 8128
rect 9377 7104 9419 7142
rect 9655 7104 9697 7142
rect 9377 7040 9385 7104
rect 9689 7040 9697 7104
rect 9377 6906 9419 7040
rect 9655 6906 9697 7040
rect 9377 6016 9697 6906
rect 9377 5952 9385 6016
rect 9449 5952 9465 6016
rect 9529 5952 9545 6016
rect 9609 5952 9625 6016
rect 9689 5952 9697 6016
rect 9377 4928 9697 5952
rect 9377 4864 9385 4928
rect 9449 4864 9465 4928
rect 9529 4864 9545 4928
rect 9609 4864 9625 4928
rect 9689 4864 9697 4928
rect 9377 3878 9697 4864
rect 9377 3840 9419 3878
rect 9655 3840 9697 3878
rect 9377 3776 9385 3840
rect 9689 3776 9697 3840
rect 9377 3642 9419 3776
rect 9655 3642 9697 3776
rect 9377 2752 9697 3642
rect 9377 2688 9385 2752
rect 9449 2688 9465 2752
rect 9529 2688 9545 2752
rect 9609 2688 9625 2752
rect 9689 2688 9697 2752
rect 9377 2128 9697 2688
<< via4 >>
rect 2672 10368 2908 10406
rect 2672 10304 2702 10368
rect 2702 10304 2718 10368
rect 2718 10304 2782 10368
rect 2782 10304 2798 10368
rect 2798 10304 2862 10368
rect 2862 10304 2878 10368
rect 2878 10304 2908 10368
rect 2672 10170 2908 10304
rect 2672 7104 2908 7142
rect 2672 7040 2702 7104
rect 2702 7040 2718 7104
rect 2718 7040 2782 7104
rect 2782 7040 2798 7104
rect 2798 7040 2862 7104
rect 2862 7040 2878 7104
rect 2878 7040 2908 7104
rect 2672 6906 2908 7040
rect 2672 3840 2908 3878
rect 2672 3776 2702 3840
rect 2702 3776 2718 3840
rect 2718 3776 2782 3840
rect 2782 3776 2798 3840
rect 2798 3776 2862 3840
rect 2862 3776 2878 3840
rect 2878 3776 2908 3840
rect 2672 3642 2908 3776
rect 4359 8736 4595 8774
rect 4359 8672 4389 8736
rect 4389 8672 4405 8736
rect 4405 8672 4469 8736
rect 4469 8672 4485 8736
rect 4485 8672 4549 8736
rect 4549 8672 4565 8736
rect 4565 8672 4595 8736
rect 4359 8538 4595 8672
rect 4359 5472 4595 5510
rect 4359 5408 4389 5472
rect 4389 5408 4405 5472
rect 4405 5408 4469 5472
rect 4469 5408 4485 5472
rect 4485 5408 4549 5472
rect 4549 5408 4565 5472
rect 4565 5408 4595 5472
rect 4359 5274 4595 5408
rect 6046 10368 6282 10406
rect 6046 10304 6076 10368
rect 6076 10304 6092 10368
rect 6092 10304 6156 10368
rect 6156 10304 6172 10368
rect 6172 10304 6236 10368
rect 6236 10304 6252 10368
rect 6252 10304 6282 10368
rect 6046 10170 6282 10304
rect 6046 7104 6282 7142
rect 6046 7040 6076 7104
rect 6076 7040 6092 7104
rect 6092 7040 6156 7104
rect 6156 7040 6172 7104
rect 6172 7040 6236 7104
rect 6236 7040 6252 7104
rect 6252 7040 6282 7104
rect 6046 6906 6282 7040
rect 6046 3840 6282 3878
rect 6046 3776 6076 3840
rect 6076 3776 6092 3840
rect 6092 3776 6156 3840
rect 6156 3776 6172 3840
rect 6172 3776 6236 3840
rect 6236 3776 6252 3840
rect 6252 3776 6282 3840
rect 6046 3642 6282 3776
rect 7732 8736 7968 8774
rect 7732 8672 7762 8736
rect 7762 8672 7778 8736
rect 7778 8672 7842 8736
rect 7842 8672 7858 8736
rect 7858 8672 7922 8736
rect 7922 8672 7938 8736
rect 7938 8672 7968 8736
rect 7732 8538 7968 8672
rect 7732 5472 7968 5510
rect 7732 5408 7762 5472
rect 7762 5408 7778 5472
rect 7778 5408 7842 5472
rect 7842 5408 7858 5472
rect 7858 5408 7922 5472
rect 7922 5408 7938 5472
rect 7938 5408 7968 5472
rect 7732 5274 7968 5408
rect 9419 10368 9655 10406
rect 9419 10304 9449 10368
rect 9449 10304 9465 10368
rect 9465 10304 9529 10368
rect 9529 10304 9545 10368
rect 9545 10304 9609 10368
rect 9609 10304 9625 10368
rect 9625 10304 9655 10368
rect 9419 10170 9655 10304
rect 9419 7104 9655 7142
rect 9419 7040 9449 7104
rect 9449 7040 9465 7104
rect 9465 7040 9529 7104
rect 9529 7040 9545 7104
rect 9545 7040 9609 7104
rect 9609 7040 9625 7104
rect 9625 7040 9655 7104
rect 9419 6906 9655 7040
rect 9419 3840 9655 3878
rect 9419 3776 9449 3840
rect 9449 3776 9465 3840
rect 9465 3776 9529 3840
rect 9529 3776 9545 3840
rect 9545 3776 9609 3840
rect 9609 3776 9625 3840
rect 9625 3776 9655 3840
rect 9419 3642 9655 3776
<< metal5 >>
rect 1104 10406 11224 10448
rect 1104 10170 2672 10406
rect 2908 10170 6046 10406
rect 6282 10170 9419 10406
rect 9655 10170 11224 10406
rect 1104 10128 11224 10170
rect 1104 8774 11224 8816
rect 1104 8538 4359 8774
rect 4595 8538 7732 8774
rect 7968 8538 11224 8774
rect 1104 8496 11224 8538
rect 1104 7142 11224 7184
rect 1104 6906 2672 7142
rect 2908 6906 6046 7142
rect 6282 6906 9419 7142
rect 9655 6906 11224 7142
rect 1104 6864 11224 6906
rect 1104 5510 11224 5552
rect 1104 5274 4359 5510
rect 4595 5274 7732 5510
rect 7968 5274 11224 5510
rect 1104 5232 11224 5274
rect 1104 3878 11224 3920
rect 1104 3642 2672 3878
rect 2908 3642 6046 3878
rect 6282 3642 9419 3878
rect 9655 3642 11224 3878
rect 1104 3600 11224 3642
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2116 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23
timestamp 1644511149
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1644511149
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95
timestamp 1644511149
transform 1 0 9844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_103
timestamp 1644511149
transform 1 0 10580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_23
timestamp 1644511149
transform 1 0 3220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_47 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1644511149
transform 1 0 6808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1644511149
transform 1 0 9016 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_98
timestamp 1644511149
transform 1 0 10120 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_106
timestamp 1644511149
transform 1 0 10856 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_17
timestamp 1644511149
transform 1 0 2668 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_25
timestamp 1644511149
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_52
timestamp 1644511149
transform 1 0 5888 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1644511149
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_95
timestamp 1644511149
transform 1 0 9844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_7
timestamp 1644511149
transform 1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_14
timestamp 1644511149
transform 1 0 2392 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_26
timestamp 1644511149
transform 1 0 3496 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_35
timestamp 1644511149
transform 1 0 4324 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1644511149
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_77
timestamp 1644511149
transform 1 0 8188 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_103
timestamp 1644511149
transform 1 0 10580 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp 1644511149
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_38
timestamp 1644511149
transform 1 0 4600 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_51
timestamp 1644511149
transform 1 0 5796 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_63
timestamp 1644511149
transform 1 0 6900 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_67
timestamp 1644511149
transform 1 0 7268 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_76
timestamp 1644511149
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_103
timestamp 1644511149
transform 1 0 10580 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_43
timestamp 1644511149
transform 1 0 5060 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1644511149
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_77
timestamp 1644511149
transform 1 0 8188 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_103
timestamp 1644511149
transform 1 0 10580 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1644511149
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_37
timestamp 1644511149
transform 1 0 4508 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_49
timestamp 1644511149
transform 1 0 5612 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_57
timestamp 1644511149
transform 1 0 6348 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1644511149
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_94
timestamp 1644511149
transform 1 0 9752 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_106
timestamp 1644511149
transform 1 0 10856 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_31
timestamp 1644511149
transform 1 0 3956 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1644511149
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_65
timestamp 1644511149
transform 1 0 7084 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_77
timestamp 1644511149
transform 1 0 8188 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_99
timestamp 1644511149
transform 1 0 10212 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_7
timestamp 1644511149
transform 1 0 1748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_19
timestamp 1644511149
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_47
timestamp 1644511149
transform 1 0 5428 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1644511149
transform 1 0 7360 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1644511149
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_95
timestamp 1644511149
transform 1 0 9844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_23
timestamp 1644511149
transform 1 0 3220 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_31
timestamp 1644511149
transform 1 0 3956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_42
timestamp 1644511149
transform 1 0 4968 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1644511149
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_65
timestamp 1644511149
transform 1 0 7084 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_75
timestamp 1644511149
transform 1 0 8004 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_103
timestamp 1644511149
transform 1 0 10580 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_11
timestamp 1644511149
transform 1 0 2116 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp 1644511149
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_49
timestamp 1644511149
transform 1 0 5612 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_55
timestamp 1644511149
transform 1 0 6164 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_76
timestamp 1644511149
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_93
timestamp 1644511149
transform 1 0 9660 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_103
timestamp 1644511149
transform 1 0 10580 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_23
timestamp 1644511149
transform 1 0 3220 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_31
timestamp 1644511149
transform 1 0 3956 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1644511149
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_65
timestamp 1644511149
transform 1 0 7084 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_89
timestamp 1644511149
transform 1 0 9292 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_101
timestamp 1644511149
transform 1 0 10396 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1644511149
transform 1 0 1748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_11
timestamp 1644511149
transform 1 0 2116 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1644511149
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_45
timestamp 1644511149
transform 1 0 5244 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_57
timestamp 1644511149
transform 1 0 6348 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1644511149
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_105
timestamp 1644511149
transform 1 0 10764 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_31
timestamp 1644511149
transform 1 0 3956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_43
timestamp 1644511149
transform 1 0 5060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_77
timestamp 1644511149
transform 1 0 8188 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_103
timestamp 1644511149
transform 1 0 10580 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_7
timestamp 1644511149
transform 1 0 1748 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1644511149
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_73
timestamp 1644511149
transform 1 0 7820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_81
timestamp 1644511149
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_94
timestamp 1644511149
transform 1 0 9752 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_101
timestamp 1644511149
transform 1 0 10396 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_24
timestamp 1644511149
transform 1 0 3312 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_48
timestamp 1644511149
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_60
timestamp 1644511149
transform 1 0 6624 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_66
timestamp 1644511149
transform 1 0 7176 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_87
timestamp 1644511149
transform 1 0 9108 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_103
timestamp 1644511149
transform 1 0 10580 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_10
timestamp 1644511149
transform 1 0 2024 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_22
timestamp 1644511149
transform 1 0 3128 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_59
timestamp 1644511149
transform 1 0 6532 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1644511149
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_103
timestamp 1644511149
transform 1 0 10580 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_7
timestamp 1644511149
transform 1 0 1748 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_20
timestamp 1644511149
transform 1 0 2944 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_35
timestamp 1644511149
transform 1 0 4324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_47
timestamp 1644511149
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_61
timestamp 1644511149
transform 1 0 6716 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_75
timestamp 1644511149
transform 1 0 8004 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_83
timestamp 1644511149
transform 1 0 8740 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_85
timestamp 1644511149
transform 1 0 8924 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_91
timestamp 1644511149
transform 1 0 9476 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_103
timestamp 1644511149
transform 1 0 10580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 11224 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 11224 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 11224 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 11224 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 11224 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 11224 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 11224 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 11224 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 11224 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 11224 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 11224 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 11224 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 11224 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 11224 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 11224 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 11224 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 11224 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 11224 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1644511149
transform 1 0 3680 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1644511149
transform 1 0 8832 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_1  _33_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2668 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _34_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _35_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _36_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 7820 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _37_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _38_
timestamp 1644511149
transform -1 0 7084 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _39_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _40_
timestamp 1644511149
transform -1 0 3220 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _41_
timestamp 1644511149
transform 1 0 4508 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _42_
timestamp 1644511149
transform -1 0 4968 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _43_
timestamp 1644511149
transform 1 0 4324 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _44_
timestamp 1644511149
transform 1 0 6164 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _45_
timestamp 1644511149
transform 1 0 5060 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _46_
timestamp 1644511149
transform 1 0 5152 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _47_
timestamp 1644511149
transform -1 0 7084 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _48_
timestamp 1644511149
transform -1 0 8004 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _49_
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _50_
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1644511149
transform 1 0 7728 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _52_
timestamp 1644511149
transform -1 0 2668 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1644511149
transform -1 0 2392 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _54_
timestamp 1644511149
transform 1 0 2208 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1644511149
transform 1 0 1840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _56_
timestamp 1644511149
transform -1 0 10580 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1644511149
transform 1 0 10120 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _58_
timestamp 1644511149
transform 1 0 4968 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1644511149
transform 1 0 4048 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _60_
timestamp 1644511149
transform -1 0 9844 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _61_
timestamp 1644511149
transform -1 0 9752 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _62_
timestamp 1644511149
transform 1 0 9108 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _63_
timestamp 1644511149
transform 1 0 7360 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _64_
timestamp 1644511149
transform -1 0 4876 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  _65_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 3220 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _66_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _67_
timestamp 1644511149
transform 1 0 5520 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _68_
timestamp 1644511149
transform -1 0 10580 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _69_
timestamp 1644511149
transform -1 0 8188 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _70_
timestamp 1644511149
transform 1 0 2116 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _71_
timestamp 1644511149
transform -1 0 3220 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _72_
timestamp 1644511149
transform 1 0 5244 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _73_
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _74_
timestamp 1644511149
transform -1 0 10580 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _75_
timestamp 1644511149
transform 1 0 7176 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _76_
timestamp 1644511149
transform 1 0 2852 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _77_
timestamp 1644511149
transform -1 0 5520 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _78_
timestamp 1644511149
transform 1 0 6256 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _79_
timestamp 1644511149
transform 1 0 8372 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _80_
timestamp 1644511149
transform -1 0 8188 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _81_
timestamp 1644511149
transform 1 0 1748 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _82_
timestamp 1644511149
transform -1 0 8464 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _83_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8464 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _84_
timestamp 1644511149
transform -1 0 5612 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _85_
timestamp 1644511149
transform 1 0 8740 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _86_
timestamp 1644511149
transform 1 0 4048 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _87_
timestamp 1644511149
transform 1 0 4048 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _88_
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _89_
timestamp 1644511149
transform 1 0 6624 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _90_
timestamp 1644511149
transform 1 0 7268 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _91_
timestamp 1644511149
transform -1 0 3220 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _92_
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _93_
timestamp 1644511149
transform 1 0 6624 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _94_
timestamp 1644511149
transform 1 0 3588 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _95_
timestamp 1644511149
transform 1 0 6624 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _96_
timestamp 1644511149
transform 1 0 6624 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _97_
timestamp 1644511149
transform -1 0 5980 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _98__17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 2024 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1644511149
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform -1 0 2944 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  input4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 10580 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  output5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10212 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1644511149
transform -1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1644511149
transform 1 0 10212 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1644511149
transform 1 0 10212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1644511149
transform 1 0 9476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1644511149
transform -1 0 9476 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1644511149
transform -1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1644511149
transform -1 0 1748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1644511149
transform 1 0 10212 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1644511149
transform 1 0 6440 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1644511149
transform -1 0 1748 0 1 9792
box -38 -48 406 592
<< labels >>
rlabel metal3 s 11529 7488 12329 7608 6 B[0]
port 0 nsew signal tristate
rlabel metal3 s 0 13608 800 13728 6 B[1]
port 1 nsew signal tristate
rlabel metal3 s 11529 10888 12329 11008 6 B[2]
port 2 nsew signal tristate
rlabel metal3 s 11529 688 12329 808 6 B[3]
port 3 nsew signal tristate
rlabel metal2 s 5814 13673 5870 14473 6 B[4]
port 4 nsew signal tristate
rlabel metal2 s 18 0 74 800 6 CompOut
port 5 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 SH
port 6 nsew signal tristate
rlabel metal5 s 1104 5232 11224 5552 6 VGND
port 7 nsew ground input
rlabel metal5 s 1104 8496 11224 8816 6 VGND
port 7 nsew ground input
rlabel metal4 s 4318 2128 4638 12016 6 VGND
port 7 nsew ground input
rlabel metal4 s 7691 2128 8011 12016 6 VGND
port 7 nsew ground input
rlabel metal5 s 1104 3600 11224 3920 6 VPWR
port 8 nsew power input
rlabel metal5 s 1104 6864 11224 7184 6 VPWR
port 8 nsew power input
rlabel metal5 s 1104 10128 11224 10448 6 VPWR
port 8 nsew power input
rlabel metal4 s 2630 2128 2950 12016 6 VPWR
port 8 nsew power input
rlabel metal4 s 6004 2128 6324 12016 6 VPWR
port 8 nsew power input
rlabel metal4 s 9377 2128 9697 12016 6 VPWR
port 8 nsew power input
rlabel metal2 s 3238 0 3294 800 6 clock
port 9 nsew signal input
rlabel metal2 s 9034 13673 9090 14473 6 dataOut[0]
port 10 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 dataOut[1]
port 11 nsew signal tristate
rlabel metal3 s 0 6808 800 6928 6 dataOut[2]
port 12 nsew signal tristate
rlabel metal2 s 12254 13673 12310 14473 6 dataOut[3]
port 13 nsew signal tristate
rlabel metal2 s 6458 0 6514 800 6 dataOut[4]
port 14 nsew signal tristate
rlabel metal3 s 0 10208 800 10328 6 nEndCnv
port 15 nsew signal tristate
rlabel metal2 s 2594 13673 2650 14473 6 nStartCnv
port 16 nsew signal input
rlabel metal3 s 11529 4088 12329 4208 6 reset
port 17 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 12329 14473
<< end >>
